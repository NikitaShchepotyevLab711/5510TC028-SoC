///////////////////////////////////////////////////////
//	File Name: test.routed.v
//	Data:      24/14/11 10:16:00
//	Program:   xcore.exe
///////////////////////////////////////////////////////
//
module test ( clk, key,  hex0,  led );
  input clk, key;
  output  [7:0] hex0;
  output  [7:0] led;
  wire \net8281<11> , \net8281<9> , \net8281<3> , \net8281<5> , \LongBus_35<10> , \LongBus_35<13> , \net8281<2> , \net8281<0> , \net8281<1> , \LongBus_35<14> , 
    \net8281<13> , \net8281<15> , \net8290<6> , \LongBus_33<9> , \LongBus_33<15> , \net8290<0> , \net8290<14> , \net8290<15> , \net8293<15> , \LongBus_30<0> , 
    \LongBus_37<4> , \net8302<11> , \LongBus_37<11> , \net8302<4> , \net8302<0> , \net8302<15> , \LongBus_37<0> , \net8305<7> , \LongBus_31<8> , \net8308<5> , 
    \net8308<7> , \net8308<1> , \net8308<15> , \net8314<11> , \net8314<7> , \net8314<15> , \LongBus_50<8> , \LongBus_50<4> , \LongBus_50<0> , \LongBus_50<15> , 
    \LongBus_11<0> , \LongBus_55<10> , \LongBus_41<14> , \LongBus_41<13> , \LongBus_41<9> , \LongBus_41<10> , \LongBus_41<11> , \LongBus_41<15> , \LongBus_40<4> , \LongBus_40<0> , 
    \LongBus_56<0> , \LongBus_56<2> , \LongBus_57<14> , \LongBus_57<12> , \LongBus_54<6> , \LongBus_54<4> , \LongBus_54<0> , \LongBus_9<8> , \LongBus_9<0> , \LongBus_10<8> , 
    \LongBus_10<0> , \LongBus_49<8> , \LongBus_49<0> , \LongBus_49<15> , \LongBus_48<9> , \LongBus_48<0> , \LongBus_48<15> , \LongBus_47<11> , \LongBus_47<4> , \LongBus_47<0> , 
    \LongBus_52<14> , \LongBus_52<0> , \LongBus_65<0> , \LongBus_63<10> , \LongBus_63<14> , \LongBus_64<4> , \LongBus_64<6> , \LongBus_64<12> , \LongBus_64<2> , \LongBus_64<0> , 
    \I3590.net78 , \I3590.net066 , \net10255<0> , \net10247<1> , \net10247<0> , \net10305<1> , \net10255<1> , \net10262<1> , \I3688.net35 , \net10244<3> , 
    \I3688.net43 , \net10244<1> , \I3688.net47 , \net10244<0> , \I3686.net35 , \net10252<3> , \I3686.net39 , \net10252<2> , \net20148<3> , \net20148<2> , 
    \GCLK_s4<0> , \GCLK_s4<2> , \GCLK_s4<3> , \IIO26.I7.net197 , \IIO26.I6.net197 , \IIO26.I5.net197 , \IIO26.I4.net197 , \IIO26.I3.net197 , \IIO26.I2.net197 , \IIO26.I1.net197 , 
    \IIO26.I0.net197 , \IIO21.I0.net0153 , \IIO21.I0.net209 , \IIO18.I7.net197 , \IIO18.I5.net197 , \IIO18.I3.net197 , \IIO18.I1.net197 , \IIO19.I7.net197 , \IIO19.I5.net197 , \IIO19.I3.net197 , 
    \IIO19.I1.net197 , \net16523<1> , \ILAB1004.I5605.net33 , \ILAB1004.Clk_int<2> , \ILAB1004.net015238 , \ILAB1004.I5366.net0119 , \LLL15_PLL1<0> , \ILAB1004.ILE1616.net01342 , \ILAB0505.I5605.net21 , \ILAB0505.Clk_int<0> , 
    \ILAB0505.I5605.net25 , \ILAB0505.Clk_int<1> , \ILAB0505.I5605.net29 , \ILAB0505.Clk_int<3> , \ILAB0505.I5605.net33 , \ILAB0505.Clk_int<2> , \ILAB0505.net27185 , \ILAB0505.net27191 , \ILAB0505.net015234 , \ILAB0505.net015238 , 
    \ILAB0505.I5366.net0122 , \net10221<0> , \net10221<1> , \ILAB0505.I5366.net0114 , \ILAB0505.net15299<3> , \ILAB0505.I5366.net0106 , \ILAB0505.net15299<1> , \ILAB0505.I5366.net0102 , \ILAB0505.net15299<0> , \ILAB0505.Clk_LAB<0> , 
    \ILAB0505.Clk_LAB<2> , \ILAB0505.Clk_LAB<3> , \ILAB0505.net24386 , \ILAB0505.net20066 , \ILAB0505.net20111 , \ILAB0505.net16016 , \net13671<1> , \ILAB0505.net38886 , \net13670<1> , \ILAB0505.net27361 , 
    \net13669<1> , \ILAB0505.net21847 , \net13670<0> , \ILAB0505.net19841 , \net14002<0> , \net13709<3> , \net13709<0> , \net13709<6> , \ILAB0505.net17914 , \ILAB0505.ILE1416.net2656 , 
    \ILAB0505.net19552 , \ILAB0505.net18067 , \ILAB0505.net19217 , \ILAB0505.ILE1413.net01345 , \ILAB0505.ILE1413.net01339 , \ILAB0505.net18364 , \ILAB0505.net19219 , \ILAB0505.ILE1413.net2656 , \net13705<1> , \net13705<3> , 
    \ILAB0505.ILE1516.net01345 , \net13705<0> , \net13705<5> , \net13705<6> , \ILAB0505.net19642 , \ILAB0505.ILE1516.net0541 , \ILAB0505.net23269 , \ILAB0505.net21262 , \ILAB0505.ILE1513.net2656 , \net14018<0> , 
    \net13659<3> , \ILAB0505.net19667 , \ILAB0505.net20409 , \net14018<1> , \ILAB0505.net19399 , \ILAB0505.ILE1412.net2656 , \ILAB0505.net24071 , \net14018<3> , \ILAB0505.net20115 , \ILAB0505.ILE1512.net2656 , 
    \net14010<0> , \ILAB0505.net22052 , \net14010<1> , \ILAB0505.net19847 , \ILAB0505.net22050 , \ILAB0505.ILE1414.net2656 , \ILAB0505.net24367 , \net14014<6> , \ILAB0505.ILE1613.net0541 , \ILAB0505.ILE1612.net01339 , 
    \net14018<6> , \net14018<5> , \net14018<4> , \ILAB0505.ILE1612.net2656 , \net13659<2> , \ILAB0505.ILE1411.net01345 , \ILAB0505.ILE1411.net2656 , \net13668<0> , \net13701<5> , \net13701<6> , 
    \net14002<6> , \ILAB0505.ILE1616.net2656 , \ILAB0505.ILE1316.net01342 , \net13713<5> , \ILAB0505.net23243 , \ILAB0505.net20972 , \ILAB0505.ILE1316.net2656 , \ILAB0505.ILE1316.net0541 , \ILAB0505.net21011 , \ILAB0505.net22226 , 
    \ILAB0505.net24682 , \ILAB0505.net20994 , \ILAB0505.ILE1313.net2656 , \ILAB0505.net21352 , \net13672<0> , \net13717<1> , \ILAB0505.net23423 , \net13717<4> , \ILAB0505.ILE1216.net2656 , \ILAB0505.ILE1312.net2656 , 
    \ILAB0505.ILE1312.net0541 , \net14022<3> , \ILAB0505.net22005 , \ILAB0505.ILE1511.net2656 , \ILAB0505.ILE1511.net0541 , \net13721<2> , \ILAB0505.ILE1611.net2656 , \ILAB0505.ILE1611.net0541 , \ILAB0505.ILE1514.net01342 , \net14010<3> , 
    \ILAB0505.ILE1514.net2656 , \ILAB0505.net24439 , \ILAB0505.net24304 , \net13659<6> , \ILAB0505.net22725 , \net14006<1> , \ILAB0505.net24257 , \ILAB0505.net22819 , \ILAB0505.net22815 , \ILAB0505.ILE1415.net2656 , 
    \ILAB0505.ILE1415.net0541 , \net14010<6> , \ILAB0505.ILE1614.net0541 , \ILAB0505.ILE1515.net2656 , \ILAB0505.ILE1314.net2656 , \ILAB0505.ILE1314.net0541 , \ILAB0505.ILE1214.net2656 , \net14026<0> , \net14026<3> , \net14026<2> , 
    \net14006<5> , \ILAB0505.ILE1615.net2656 , \ILAB0505.net24302 , \ILAB0505.ILE1315.net2656 , \ILAB0505.ILE1610.net0560 , \net14026<6> , \ILAB0505.ILE1610.net2656 , \ILAB0505.ILE1610.net0541 , \ILAB0505.net24435 , \ILAB0505.ILE1215.net0560 , 
    \ILAB0505.ILE1215.net2656 , \ILAB0505.ILE1115.net2656 , \ILAB0605.I5366.net64 , \ILAB0605.I5366.net66 , \ILAB0605.I5366.net68 , \net10229<0> , \net10229<1> , \ILAB0605.I5366.net0114 , \ILAB0605.net15299<3> , \ILAB0605.I5366.net0106 , 
    \ILAB0605.net15299<1> , \ILAB0605.I5366.net0102 , \ILAB0605.net15299<0> , \ILAB0605.Clk_LAB<0> , \ILAB0605.Clk_LAB<2> , \ILAB0605.Clk_LAB<3> , \ILAB0605.net21911 , \ILAB0605.net25852 , \ILAB0605.net17077 , \ILAB0605.net16339 , 
    \ILAB0605.net15439 , \ILAB0605.net16807 , \ILAB0605.net16511 , \ILAB0605.net18112 , \ILAB0605.net16672 , \net13981<0> , \ILAB0605.net19796 , \net14047<1> , \net14047<2> , \net14047<3> , 
    \ILAB0605.ILE0516.net01339 , \ILAB0605.ILE0516.net01342 , \net14047<0> , \net14047<6> , \ILAB0605.net19057 , \ILAB0605.net17014 , \ILAB0605.net18859 , \ILAB0605.ILE0516.net2656 , \net13982<0> , \ILAB0605.net19256 , 
    \net14051<3> , \ILAB0605.ILE0416.net0562 , \net14051<6> , \ILAB0605.ILE0416.net2656 , \ILAB0605.net19984 , \ILAB0605.net19352 , \ILAB0605.net20362 , \ILAB0605.ILE0513.net0562 , \ILAB0605.net23917 , \ILAB0605.net25519 , 
    \ILAB0605.net18319 , \ILAB0605.net19354 , \ILAB0605.ILE0513.net2656 , \ILAB0605.net18499 , \ILAB0605.net18949 , \net14043<1> , \ILAB0605.net23964 , \net14043<2> , \ILAB0605.ILE0616.net01342 , \net14043<0> , 
    \net14043<4> , \ILAB0605.ILE0616.net2656 , \ILAB0605.net19031 , \ILAB0605.ILE0412.net0562 , \ILAB0605.ILE0412.net01339 , \ILAB0605.ILE0412.net2656 , \ILAB0605.net23936 , \ILAB0605.net20364 , \ILAB0605.ILE0512.net2656 , \ILAB0605.net19121 , 
    \ILAB0605.net22144 , \ILAB0605.ILE0414.net0562 , \ILAB0605.net19262 , \ILAB0605.net19804 , \ILAB0605.ILE0414.net2656 , \ILAB0605.net19346 , \ILAB0605.net21461 , \ILAB0605.net21442 , \ILAB0605.net19706 , \ILAB0605.net24097 , 
    \ILAB0605.ILE0613.net2656 , \ILAB0605.ILE0613.net0541 , \ILAB0605.net21444 , \ILAB0605.ILE0612.net0541 , \ILAB0605.ILE0514.net0558 , \ILAB0605.ILE0514.net2656 , \ILAB0605.net21469 , \ILAB0605.ILE0411.net0562 , \ILAB0605.net19892 , \ILAB0605.net21467 , 
    \ILAB0605.net20389 , \ILAB0605.ILE0411.net2656 , \ILAB0605.net23919 , \ILAB0605.ILE0511.net2656 , \ILAB0605.ILE0511.net0541 , \ILAB0605.ILE0611.net01345 , \ILAB0605.ILE0611.net2656 , \ILAB0605.ILE0711.net01345 , \ILAB0605.ILE0711.net2656 , \net14063<1> , 
    \net14063<3> , \ILAB0605.ILE0116.net0562 , \ILAB0605.ILE0116.net0558 , \net14063<0> , \net14063<6> , \ILAB0605.net21892 , \ILAB0605.ILE0116.net2656 , \ILAB0605.net23197 , \ILAB0605.ILE0112.net0562 , \ILAB0605.net21894 , 
    \ILAB0605.ILE0112.net2656 , \ILAB0605.net23756 , \net14059<1> , \net14059<2> , \net14059<6> , \ILAB0605.ILE0216.net2656 , \ILAB0605.net22099 , \ILAB0605.ILE0614.net2656 , \ILAB0605.ILE0614.net0541 , \ILAB0605.ILE0113.net01342 , 
    \ILAB0605.net23177 , \ILAB0605.net23085 , \ILAB0605.ILE0113.net2656 , \ILAB0605.ILE0113.net0541 , \ILAB0605.net22316 , \ILAB0605.ILE0212.net01342 , \ILAB0605.net23306 , \ILAB0605.net22299 , \ILAB0605.ILE0212.net2656 , \ILAB0605.ILE0212.net0541 , 
    \ILAB0605.net22367 , \ILAB0605.net22459 , \ILAB0605.net22455 , \ILAB0605.ILE0415.net0541 , \ILAB0605.ILE0515.net2656 , \ILAB0605.ILE0515.net0541 , \net14055<1> , \ILAB0605.net24819 , \net14055<3> , \ILAB0605.ILE0316.net0560 , 
    \net14055<0> , \net14055<5> , \net14055<6> , \ILAB0605.ILE0316.net2656 , \ILAB0605.ILE0213.net0541 , \ILAB0605.net24909 , \ILAB0605.net24926 , \ILAB0605.net25897 , \ILAB0605.net23153 , \ILAB0605.net26100 , 
    \ILAB0605.ILE0313.net2656 , \ILAB0605.ILE0313.net0541 , \ILAB0605.ILE0111.net01345 , \ILAB0605.ILE0111.net0560 , \ILAB0605.ILE0111.net2656 , \ILAB0605.ILE0211.net0562 , \ILAB0605.ILE0211.net2656 , \ILAB0605.net25899 , \ILAB0605.ILE0311.net2656 , \ILAB0605.net23629 , 
    \ILAB0605.net23807 , \ILAB0605.ILE0114.net2656 , \ILAB0605.ILE0214.net01345 , \ILAB0605.ILE0214.net2656 , \ILAB0605.ILE0314.net2656 , \ILAB0605.net23942 , \ILAB0605.net23897 , \ILAB0605.ILE0410.net2656 , \ILAB0605.ILE0510.net2656 , \ILAB0605.ILE0510.net0541 , 
    \ILAB0605.ILE0615.net2656 , \ILAB0605.ILE0115.net01342 , \ILAB0605.net24842 , \ILAB0605.net24615 , \ILAB0605.ILE0115.net2656 , \ILAB0605.ILE0215.net2656 , \ILAB0605.ILE0215.net0541 , \ILAB0605.ILE0315.net2656 , \ILAB0605.ILE0312.net0558 , \ILAB0605.ILE0312.net2656 , 
    \ILAB0605.ILE0110.net2656 , \ILAB0605.ILE0310.net2656 , \ILAB0605.ILE0310.net0541 , \ILAB0605.ILE0413.net2656 , \ILAB0605.ILE0413.net0541 , \ILAB0506.I5605.net21 , \ILAB0506.Clk_int<0> , \ILAB0506.I5605.net25 , \ILAB0506.Clk_int<1> , \ILAB0506.I5605.net29 , 
    \ILAB0506.Clk_int<3> , \ILAB0506.I5605.net33 , \ILAB0506.Clk_int<2> , \ILAB0506.net027160 , \ILAB0506.net027166 , \ILAB0506.net27188 , \ILAB0506.net27128 , \ILAB0506.I5366.net0119 , \ILAB0506.I5366.net0110 , \ILAB0506.net15299<2> , 
    \ILAB0506.I5366.net0106 , \ILAB0506.net15299<1> , \ILAB0506.I5366.net0102 , \ILAB0506.net15299<0> , \ILAB0506.Clk_LAB<1> , \ILAB0506.Clk_LAB<2> , \ILAB0506.Clk_LAB<3> , \ILAB0506.net15881 , \ILAB0506.net25376 , \ILAB0506.net15476 , 
    \ILAB0506.net20561 , \net14730<1> , \ILAB0506.net27283 , \net14735<1> , \ILAB0506.net27289 , \net14732<1> , \ILAB0506.net27297 , \net14738<1> , \ILAB0506.net27303 , \net14736<1> , 
    \ILAB0506.net27339 , \net15095<1> , \ILAB0506.net19597 , \net15111<3> , \net15111<1> , \ILAB0506.ILE1603.net01345 , \ILAB0506.net15458 , \net15111<6> , \ILAB0506.net15484 , \ILAB0506.net15459 , 
    \net15111<4> , \ILAB0506.ILE1603.net2656 , \ILAB0506.net15521 , \ILAB0506.net20839 , \ILAB0506.ILE1201.net0560 , \ILAB0506.ILE1201.net0541 , \ILAB0506.net20029 , \ILAB0506.net17726 , \net15103<1> , \ILAB0506.net20857 , 
    \ILAB0506.ILE1605.net0560 , \ILAB0506.ILE1605.net0558 , \ILAB0506.net25067 , \ILAB0506.net15908 , \net15107<1> , \ILAB0506.net25382 , \ILAB0506.net25384 , \ILAB0506.ILE1504.net0541 , \ILAB0506.net18049 , \ILAB0506.net18697 , 
    \ILAB0506.net25807 , \ILAB0506.ILE1101.net01339 , \ILAB0506.net16584 , \net14802<1> , \ILAB0506.net17149 , \ILAB0506.net18922 , \ILAB0506.ILE1503.net01345 , \ILAB0506.ILE1503.net0560 , \ILAB0506.net20858 , \ILAB0506.ILE1503.net2656 , 
    \net15099<3> , \ILAB0506.ILE1606.net0562 , \ILAB0506.ILE1606.net0558 , \net15099<6> , \net15099<4> , \ILAB0506.ILE1606.net2656 , \ILAB0506.net18311 , \ILAB0506.net22549 , \ILAB0506.net19984 , \ILAB0506.net19354 , 
    \ILAB0506.net18499 , \ILAB0506.net21694 , \ILAB0506.net21692 , \ILAB0506.net19687 , \ILAB0506.net23539 , \ILAB0506.net23494 , \ILAB0506.net18904 , \ILAB0506.net18967 , \ILAB0506.net18986 , \ILAB0506.net25312 , 
    \ILAB0506.net21690 , \ILAB0506.ILE0912.net2656 , \ILAB0506.ILE0912.net0541 , \ILAB0506.net19031 , \ILAB0506.net19939 , \ILAB0506.net19082 , \net14773<6> , \ILAB0506.net19084 , \ILAB0506.net19014 , \ILAB0506.ILE0412.net2656 , 
    \ILAB0506.ILE0512.net01345 , \ILAB0506.ILE0512.net2656 , \ILAB0506.net25493 , \ILAB0506.net23537 , \ILAB0506.ILE0914.net2656 , \ILAB0506.net22414 , \ILAB0506.net22144 , \ILAB0506.net26078 , \ILAB0506.net19804 , \ILAB0506.ILE0414.net2656 , 
    \net14734<0> , \net14794<1> , \ILAB0506.ILE0716.net01345 , \ILAB0506.net19346 , \ILAB0506.net21442 , \ILAB0506.ILE0613.net0562 , \ILAB0506.net21443 , \ILAB0506.net21424 , \ILAB0506.ILE0613.net2656 , \ILAB0506.net24116 , 
    \ILAB0506.net24098 , \ILAB0506.ILE0612.net2656 , \ILAB0506.ILE0514.net2656 , \ILAB0506.ILE0514.net0541 , \ILAB0506.net21514 , \ILAB0506.net21469 , \ILAB0506.net20387 , \ILAB0506.ILE0411.net01339 , \ILAB0506.net20389 , \ILAB0506.ILE0411.net2656 , 
    \ILAB0506.ILE0712.net01345 , \ILAB0506.ILE0712.net2656 , \ILAB0506.net19976 , \ILAB0506.net19959 , \ILAB0506.ILE0713.net2656 , \ILAB0506.net20021 , \ILAB0506.net20812 , \ILAB0506.net26303 , \ILAB0506.net26302 , \ILAB0506.net20003 , 
    \ILAB0506.ILE1403.net2656 , \ILAB0506.ILE0511.net2656 , \ILAB0506.ILE1301.net01339 , \net15119<0> , \ILAB0506.ILE1301.net2656 , \net15119<3> , \net15119<1> , \ILAB0506.ILE1601.net01342 , \net15119<5> , \ILAB0506.ILE1601.net0541 , 
    \ILAB0506.net20814 , \ILAB0506.ILE1401.net2656 , \ILAB0506.ILE1401.net0541 , \ILAB0506.ILE1501.net2656 , \ILAB0506.net24682 , \ILAB0506.net21416 , \ILAB0506.net22676 , \ILAB0506.net22657 , \ILAB0506.ILE1013.net01345 , \ILAB0506.net24862 , 
    \ILAB0506.ILE1013.net2656 , \ILAB0506.ILE0611.net2656 , \ILAB0506.ILE0611.net0541 , \ILAB0506.net21759 , \ILAB0506.ILE1113.net01339 , \ILAB0506.net24952 , \ILAB0506.net21534 , \ILAB0506.ILE1113.net2656 , \ILAB0506.ILE1012.net2656 , \ILAB0506.ILE1012.net0541 , 
    \net14778<1> , \ILAB0506.ILE1112.net2656 , \ILAB0506.net22099 , \ILAB0506.net22189 , \ILAB0506.ILE0614.net2656 , \ILAB0506.ILE0614.net0541 , \ILAB0506.ILE0915.net2656 , \ILAB0506.ILE0415.net0562 , \ILAB0506.ILE0415.net2656 , \ILAB0506.ILE0714.net2656 , 
    \ILAB0506.ILE0714.net0541 , \ILAB0506.ILE0515.net0562 , \ILAB0506.ILE0515.net0558 , \ILAB0506.ILE0515.net2656 , \ILAB0506.net24819 , \net14810<0> , \ILAB0506.ILE0813.net01345 , \ILAB0506.ILE0813.net2656 , \ILAB0506.net23396 , \ILAB0506.net23153 , 
    \ILAB0506.ILE0313.net2656 , \net14777<1> , \ILAB0506.ILE0311.net2656 , \ILAB0506.ILE1014.net2656 , \ILAB0506.ILE1014.net0541 , \ILAB0506.ILE1114.net2656 , \net14765<1> , \ILAB0506.ILE0314.net2656 , \ILAB0506.ILE0615.net2656 , \ILAB0506.ILE0312.net2656 , 
    \ILAB0506.ILE0312.net0541 , \ILAB0506.ILE1405.net2656 , \ILAB0506.ILE1604.net0560 , \net15107<6> , \net15107<5> , \ILAB0506.ILE1604.net2656 , \ILAB0506.ILE1604.net0541 , \ILAB0506.ILE0913.net0562 , \ILAB0506.ILE0913.net2656 , \ILAB0506.ILE1404.net2656 , 
    \ILAB0506.ILE1404.net0541 , \ILAB0506.ILE0413.net0541 , \ILAB0506.net26554 , \net15115<0> , \ILAB0506.net26509 , \net15115<1> , \ILAB0506.ILE1402.net2656 , \ILAB0506.ILE1502.net2656 , \ILAB0506.ILE1602.net0541 , \ILAB0506.ILE1302.net0558 , 
    \ILAB0506.ILE1302.net01342 , \ILAB0506.ILE1302.net2656 , \ILAB0506.ILE1202.net0541 , \ILAB0706.I5366.net64 , \ILAB0706.I5366.net70 , \ILAB0706.I5366.net0114 , \ILAB0706.net15299<3> , \ILAB0706.I5366.net0110 , \ILAB0706.net15299<2> , \ILAB0706.Clk_LAB<0> , 
    \ILAB0706.Clk_LAB<1> , \ILAB0706.net22271 , \ILAB0706.net38763 , \ILAB0706.net23666 , \ILAB0706.net38388 , \ILAB0706.net21911 , \ILAB0706.net38625 , \net14936<1> , \net14916<6> , \net14924<2> , 
    \ILAB0706.net22320 , \net14920<6> , \ILAB0706.ILE0113.net0541 , \net14912<6> , \net14928<0> , \net14928<1> , \net14916<3> , \net14916<4> , \net14916<1> , \ILAB0706.ILE0114.net0541 , 
    \ILAB0706.ILE0115.net0541 , \net14932<4> , \net14932<5> , \net14932<0> , \ILAB0606.I5605.net21 , \ILAB0606.Clk_int<0> , \ILAB0606.I5605.net25 , \ILAB0606.Clk_int<1> , \ILAB0606.I5605.net33 , \ILAB0606.Clk_int<2> , 
    \ILAB0606.net27185 , \ILAB0606.net27191 , \ILAB0606.net015238 , \ILAB0606.I5366.net0122 , \ILAB0606.I5366.net0119 , \ILAB0606.I5366.net0106 , \ILAB0606.net15299<1> , \ILAB0606.Clk_LAB<2> , \ILAB0606.net24386 , \ILAB0606.net20066 , 
    \ILAB0606.net22766 , \ILAB0606.net20111 , \ILAB0606.net21641 , \ILAB0606.net38760 , \net15030<1> , \ILAB0606.net27307 , \ILAB0606.net22946 , \ILAB0606.net19751 , \net15029<1> , \ILAB0606.net27361 , 
    \net15028<1> , \ILAB0606.net27381 , \ILAB0606.net39819 , \ILAB0606.net15349 , \ILAB0606.net25852 , \ILAB0606.net17528 , \ILAB0606.net16132 , \ILAB0606.net17644 , \ILAB0606.net15566 , \ILAB0606.net26231 , 
    \ILAB0606.net16114 , \ILAB0606.net25022 , \ILAB0606.net26212 , \ILAB0606.net20182 , \ILAB0606.net15548 , \ILAB0606.net26213 , \ILAB0606.ILE0404.net2656 , \ILAB0606.net15799 , \ILAB0606.net16020 , \ILAB0606.ILE1609.net0562 , 
    \ILAB0606.ILE1609.net0558 , \ILAB0606.net26797 , \ILAB0606.net23557 , \ILAB0606.net23576 , \ILAB0606.net26798 , \ILAB0606.ILE0304.net2656 , \ILAB0606.ILE0304.net0541 , \ILAB0606.net16241 , \ILAB0606.net18049 , \ILAB0606.net18092 , 
    \ILAB0606.net17122 , \ILAB0606.net21866 , \ILAB0606.net16222 , \ILAB0606.net18047 , \ILAB0606.net16249 , \ILAB0606.net18094 , \ILAB0606.ILE1309.net2656 , \ILAB0606.ILE1309.net0541 , \ILAB0606.net16292 , \ILAB0606.net16294 , 
    \ILAB0606.ILE1209.net2656 , \ILAB0606.net24772 , \ILAB0606.net16358 , \ILAB0606.ILE1109.net2656 , \ILAB0606.net17257 , \ILAB0606.net16403 , \ILAB0606.net25249 , \net15022<6> , \ILAB0606.net16717 , \ILAB0606.net17867 , 
    \ILAB0606.ILE0101.net2656 , \ILAB0606.net20137 , \ILAB0606.ILE0107.net01342 , \ILAB0606.ILE0107.net2656 , \ILAB0606.net20227 , \ILAB0606.net23827 , \ILAB0606.ILE0207.net2656 , \ILAB0606.net16943 , \ILAB0606.net16944 , \ILAB0606.ILE0201.net2656 , 
    \ILAB0606.net17059 , \ILAB0606.ILE0106.net01342 , \ILAB0606.net22928 , \ILAB0606.net26707 , \net15022<5> , \ILAB0606.net17552 , \ILAB0606.ILE0106.net2656 , \ILAB0606.ILE0106.net0541 , \ILAB0606.net18589 , \ILAB0606.net23334 , 
    \ILAB0606.net23351 , \ILAB0606.ILE0306.net2656 , \ILAB0606.ILE0306.net0541 , \ILAB0606.net17685 , \ILAB0606.net17687 , \ILAB0606.net17689 , \ILAB0606.ILE0405.net01342 , \ILAB0606.ILE0405.net0541 , \ILAB0606.ILE0301.net0562 , \ILAB0606.ILE0301.net01342 , 
    \ILAB0606.net17843 , \ILAB0606.net20524 , \ILAB0606.net20745 , \ILAB0606.ILE0301.net2656 , \ILAB0606.net19841 , \net15068<2> , \net15068<0> , \ILAB0606.net19372 , \ILAB0606.ILE0406.net2656 , \ILAB0606.net18356 , 
    \ILAB0606.net19373 , \ILAB0606.net18338 , \ILAB0606.ILE1413.net2656 , \ILAB0606.net26752 , \ILAB0606.ILE0206.net2656 , \ILAB0606.net22682 , \ILAB0606.net18994 , \ILAB0606.net21784 , \ILAB0606.ILE0506.net01339 , \ILAB0606.ILE0506.net2656 , 
    \ILAB0606.net22046 , \net15064<0> , \ILAB0606.net23539 , \ILAB0606.net23449 , \ILAB0606.net21262 , \ILAB0606.net19643 , \ILAB0606.ILE1513.net2656 , \ILAB0606.net19397 , \ILAB0606.net19399 , \ILAB0606.ILE1412.net2656 , 
    \ILAB0606.ILE1512.net2656 , \ILAB0606.net23357 , \ILAB0606.ILE0105.net0541 , \ILAB0606.net22772 , \ILAB0606.net22054 , \ILAB0606.ILE1414.net2656 , \ILAB0606.ILE1414.net0541 , \ILAB0606.net20092 , \ILAB0606.ILE1613.net2656 , \ILAB0606.ILE1613.net0541 , 
    \ILAB0606.ILE1612.net2656 , \ILAB0606.net20632 , \ILAB0606.net26258 , \ILAB0606.net20162 , \ILAB0606.ILE0503.net2656 , \ILAB0606.net20741 , \ILAB0606.net26214 , \ILAB0606.ILE0403.net01339 , \ILAB0606.net20723 , \ILAB0606.ILE0403.net2656 , 
    \ILAB0606.ILE0403.net0541 , \ILAB0606.ILE0204.net2656 , \net15018<2> , \ILAB0606.ILE1411.net01339 , \ILAB0606.ILE1411.net2656 , \ILAB0606.ILE0601.net01342 , \ILAB0606.ILE0601.net2656 , \ILAB0606.ILE0501.net2656 , \ILAB0606.ILE0501.net0541 , \ILAB0606.ILE0401.net0541 , 
    \net15072<0> , \ILAB0606.net21011 , \ILAB0606.net22226 , \ILAB0606.net21219 , \ILAB0606.net21218 , \ILAB0606.net24682 , \ILAB0606.net20993 , \ILAB0606.ILE1313.net2656 , \ILAB0606.net22586 , \ILAB0606.net22567 , 
    \ILAB0606.net21354 , \ILAB0606.ILE1213.net01345 , \ILAB0606.ILE1213.net0558 , \ILAB0606.net21083 , \ILAB0606.net21109 , \ILAB0606.ILE1213.net2656 , \ILAB0606.net21242 , \ILAB0606.ILE1312.net2656 , \ILAB0606.ILE1312.net0541 , \ILAB0606.ILE1511.net2656 , 
    \ILAB0606.ILE0205.net0558 , \ILAB0606.ILE0205.net01342 , \ILAB0606.ILE0205.net2656 , \ILAB0606.net24728 , \ILAB0606.ILE1212.net0541 , \ILAB0606.net21686 , \ILAB0606.net24862 , \ILAB0606.ILE1013.net0541 , \ILAB0606.net21551 , \ILAB0606.net23017 , 
    \ILAB0606.net21758 , \ILAB0606.net23018 , \ILAB0606.ILE1016.net01339 , \ILAB0606.ILE1112.net2656 , \ILAB0606.net23199 , \ILAB0606.ILE1611.net0541 , \ILAB0606.ILE1514.net2656 , \ILAB0606.net24684 , \ILAB0606.ILE1311.net2656 , \ILAB0606.net23783 , 
    \ILAB0606.net24729 , \ILAB0606.ILE1211.net2656 , \ILAB0606.net23040 , \ILAB0606.ILE1415.net0541 , \ILAB0606.ILE1614.net2656 , \ILAB0606.ILE1614.net0541 , \ILAB0606.ILE1515.net01345 , \ILAB0606.ILE1515.net0541 , \ILAB0606.ILE0103.net01339 , \ILAB0606.net23582 , 
    \ILAB0606.ILE0103.net2656 , \ILAB0606.ILE0104.net2656 , \ILAB0606.ILE1111.net0562 , \ILAB0606.ILE1111.net2656 , \ILAB0606.net23377 , \ILAB0606.net24909 , \ILAB0606.ILE0305.net2656 , \ILAB0606.net25898 , \ILAB0606.ILE1214.net2656 , \ILAB0606.ILE1014.net2656 , 
    \ILAB0606.ILE1114.net01345 , \ILAB0606.ILE1114.net2656 , \ILAB0606.ILE1114.net0541 , \ILAB0606.net26799 , \ILAB0606.ILE0303.net2656 , \ILAB0606.ILE0203.net2656 , \ILAB0606.net24077 , \ILAB0606.ILE1410.net01345 , \ILAB0606.ILE1410.net01339 , \ILAB0606.net24032 , 
    \ILAB0606.net24392 , \ILAB0606.net24034 , \ILAB0606.net24079 , \ILAB0606.net24075 , \ILAB0606.ILE1410.net2656 , \ILAB0606.net24390 , \ILAB0606.ILE1615.net2656 , \ILAB0606.ILE1615.net0541 , \ILAB0606.ILE1610.net0560 , \ILAB0606.ILE1310.net2656 , 
    \ILAB0606.ILE1310.net0541 , \ILAB0606.ILE1210.net2656 , \ILAB0606.ILE1110.net2656 , \ILAB0606.ILE0504.net2656 , \ILAB0606.ILE0505.net2656 , \ILAB0606.net26464 , \ILAB0606.net26237 , \net15022<1> , \ILAB0606.ILE0402.net2656 , \ILAB0606.ILE0402.net0541 , 
    \ILAB0606.ILE0502.net01339 , \ILAB0606.ILE0502.net2656 , \ILAB0606.net26822 , \ILAB0606.ILE0102.net2656 , \ILAB0606.ILE0202.net2656 , \ILAB0606.ILE0302.net2656 , \ILAB0406.net24386 , \ILAB0406.net20066 , \ILAB0406.net38760 , \ILAB0406.net37986 , 
    \ILAB0507.net39618 , \ILAB0507.ILE1101.net01339 , \ILAB0507.ILE0701.net01339 , \ILAB0507.ILE0601.net01339 , \ILAB0507.ILE0501.net01339 , \ILAB0607.ILE1101.net01339 , \IIO30.I7.net0151 , \IIO30.I7.net0153 , \IIO30.I7.net209 ,
    GND, VDD;
  assign GND = 1'b0;
  assign VDD = 1'b1;

  //initial $sdf_annotate("C:/Users/Admin-PC/Desktop/xcad_projects/test/prj/test.STA.reports/test.routed.sdf");

  xci2_ib XC_BUF_clk ( .a(clk), .x(\IIO30.I7.net209 ));
  xci2_ib XC_BUF_key ( .a(key), .x(\IIO21.I0.net209 ));
  xci2_ob \XC_BUF_hex0[0]  ( .a(\IIO26.I0.net197 ), .x(hex0[0]));
  xci2_ob \XC_BUF_hex0[1]  ( .a(\IIO26.I1.net197 ), .x(hex0[1]));
  xci2_ob \XC_BUF_hex0[2]  ( .a(\IIO26.I2.net197 ), .x(hex0[2]));
  xci2_ob \XC_BUF_hex0[3]  ( .a(\IIO26.I3.net197 ), .x(hex0[3]));
  xci2_ob \XC_BUF_hex0[4]  ( .a(\IIO26.I4.net197 ), .x(hex0[4]));
  xci2_ob \XC_BUF_hex0[5]  ( .a(\IIO26.I5.net197 ), .x(hex0[5]));
  xci2_ob \XC_BUF_hex0[6]  ( .a(\IIO26.I6.net197 ), .x(hex0[6]));
  xci2_ob \XC_BUF_hex0[7]  ( .a(\IIO26.I7.net197 ), .x(hex0[7]));
  xci2_ob \XC_BUF_led[0]  ( .a(\IIO19.I1.net197 ), .x(led[0]));
  xci2_ob \XC_BUF_led[1]  ( .a(\IIO19.I3.net197 ), .x(led[1]));
  xci2_ob \XC_BUF_led[2]  ( .a(\IIO19.I5.net197 ), .x(led[2]));
  xci2_ob \XC_BUF_led[3]  ( .a(\IIO19.I7.net197 ), .x(led[3]));
  xci2_ob \XC_BUF_led[4]  ( .a(\IIO18.I1.net197 ), .x(led[4]));
  xci2_ob \XC_BUF_led[5]  ( .a(\IIO18.I3.net197 ), .x(led[5]));
  xci2_ob \XC_BUF_led[6]  ( .a(\IIO18.I5.net197 ), .x(led[6]));
  xci2_ob \XC_BUF_led[7]  ( .a(\IIO18.I7.net197 ), .x(led[7]));
  xci2_nor2 _143_ ( .a(\net15111<4> ), .b(\ILAB0606.ILE0103.net01339 ), .y(\ILAB0606.ILE0103.net2656 ));
  xci2_and3fft _144_ ( .a(\ILAB0506.net20858 ), .b(\ILAB0605.net24842 ), .c(\net14063<3> ), .y(\ILAB0606.ILE0101.net2656 ));
  xci2_nor2 _145_ ( .a(\ILAB0505.Clk_LAB<2> ), .b(\net14018<5> ), .y(\ILAB0505.ILE1613.net0541 ));
  xci2_and3fft _146_ ( .a(\ILAB0505.net22052 ), .b(\ILAB0505.net19847 ), .c(\ILAB0505.Clk_LAB<0> ), .y(\ILAB0505.ILE1414.net2656 ));
  xci2_nor2 _147_ ( .a(\ILAB0605.ILE0414.net0562 ), .b(\ILAB0605.net19352 ), .y(\ILAB0605.ILE0414.net2656 ));
  xci2_and3fft _148_ ( .a(\net14055<0> ), .b(\ILAB0605.net26100 ), .c(\net14010<6> ), .y(\ILAB0605.ILE0314.net2656 ));
  xci2_and3 _149_ ( .a(\net14063<0> ), .b(\net14010<1> ), .c(\ILAB0605.net23197 ), .y(\ILAB0605.ILE0114.net2656 ));
  xci2_and2 _150_ ( .a(\ILAB0605.net23919 ), .b(\ILAB0605.net18499 ), .y(\ILAB0605.ILE0511.net2656 ));
  xci2_and2 _150__1 ( .a(\ILAB0605.net23919 ), .b(\ILAB0605.net18499 ), .y(\ILAB0605.ILE0511.net0541 ));
  xci2_and2 _151_ ( .a(\ILAB0505.net22725 ), .b(\ILAB0506.ILE1301.net01339 ), .y(\ILAB0506.ILE1301.net2656 ));
  xci2_nor2 _152_ ( .a(\net15107<5> ), .b(\net15107<1> ), .y(\ILAB0606.ILE0104.net2656 ));
  xci2_and3 _153_ ( .a(\net14059<2> ), .b(\net15119<5> ), .c(\ILAB0606.net16717 ), .y(\ILAB0606.ILE0201.net2656 ));
  xci2_nor2 _154_ ( .a(\net15099<3> ), .b(\net15099<6> ), .y(\ILAB0606.ILE0206.net2656 ));
  xci2_and3fft _155_ ( .a(\ILAB0606.net26237 ), .b(\net15107<6> ), .c(\ILAB0606.net26752 ), .y(\ILAB0606.ILE0204.net2656 ));
  xci2_and2 _156_ ( .a(\ILAB0505.net21262 ), .b(\ILAB0505.net24257 ), .y(\ILAB0505.ILE1614.net0541 ));
  xci2_and3 _157_ ( .a(\ILAB0605.net22459 ), .b(\ILAB0605.net23153 ), .c(\ILAB0605.Clk_LAB<3> ), .y(\ILAB0605.ILE0315.net2656 ));
  xci2_and3 _158_ ( .a(\ILAB0606.net16944 ), .b(\net14059<6> ), .c(\ILAB0606.net26822 ), .y(\ILAB0606.ILE0202.net2656 ));
  xci2_and2 _159_ ( .a(\net14063<1> ), .b(\net15115<1> ), .y(\ILAB0606.ILE0102.net2656 ));
  xci2_nand3ftt _160_ ( .a(\ILAB0606.ILE0301.net0562 ), .b(\ILAB0606.ILE0301.net01342 ), .c(\net15119<3> ), .y(\ILAB0606.ILE0301.net2656 ));
  xci2_and3fft _161_ ( .a(\ILAB0606.net17843 ), .b(\net14055<1> ), .c(\ILAB0606.net20745 ), .y(\ILAB0606.ILE0302.net2656 ));
  xci2_and3fft _162_ ( .a(\ILAB0605.ILE0214.net01345 ), .b(\ILAB0605.net19804 ), .c(\ILAB0605.net20364 ), .y(\ILAB0605.ILE0214.net2656 ));
  xci2_and3fft _163_ ( .a(\net14051<3> ), .b(\ILAB0506.net15458 ), .c(\ILAB0606.net16943 ), .y(\ILAB0606.ILE0203.net2656 ));
  xci2_nor3 _164_ ( .a(\ILAB0605.ILE0416.net0562 ), .b(\net14055<5> ), .c(\ILAB0605.net22455 ), .y(\ILAB0605.ILE0416.net2656 ));
  xci2_or2 _165_ ( .a(\ILAB0506.net26303 ), .b(\ILAB0506.net26509 ), .y(\ILAB0506.ILE1602.net0541 ));
  xci2_and3fft _166_ ( .a(\ILAB0605.net19352 ), .b(\ILAB0605.Clk_LAB<0> ), .c(\ILAB0605.net24819 ), .y(\ILAB0605.ILE0415.net0541 ));
  xci2_nand3ftt _167_ ( .a(\ILAB0505.net22052 ), .b(\ILAB0505.ILE1514.net01342 ), .c(\ILAB0505.net21262 ), .y(\ILAB0505.ILE1514.net2656 ));
  xci2_and3fft _168_ ( .a(\ILAB0605.net19262 ), .b(\ILAB0605.net17014 ), .c(\net14063<6> ), .y(\ILAB0605.ILE0216.net2656 ));
  xci2_and3 _169_ ( .a(\net14002<6> ), .b(\ILAB0605.ILE0316.net0560 ), .c(\ILAB0605.net18859 ), .y(\ILAB0605.ILE0316.net2656 ));
  xci2_nand3 _170_ ( .a(\ILAB0606.net26799 ), .b(\ILAB0606.net17689 ), .c(\net14055<6> ), .y(\ILAB0606.ILE0303.net2656 ));
  xci2_and2ft _171_ ( .a(\ILAB0506.net15908 ), .b(\ILAB0506.ILE1605.net0558 ), .y(\ILAB0506.ILE1405.net2656 ));
  xci2_and3ftt _172_ ( .a(\net15095<1> ), .b(\ILAB0606.net23582 ), .c(\ILAB0606.ILE0107.net01342 ), .y(\ILAB0606.ILE0107.net2656 ));
  xci2_xnor2ft _173_ ( .a(\ILAB0606.net23827 ), .b(\ILAB0606.net22928 ), .y(\ILAB0606.ILE0105.net0541 ));
  xci2_and3 _174_ ( .a(\ILAB0506.ILE1606.net0562 ), .b(\net15111<6> ), .c(\ILAB0506.ILE1606.net0558 ), .y(\ILAB0506.ILE1606.net2656 ));
  xci2_aoi21 _175_ ( .a(\ILAB0606.net23827 ), .b(\ILAB0606.ILE0205.net01342 ), .c(\ILAB0606.ILE0205.net0558 ), .y(\ILAB0606.ILE0205.net2656 ));
  xci2_and3 _176_ ( .a(\ILAB0606.net20227 ), .b(\ILAB0606.net22928 ), .c(\ILAB0606.net26797 ), .y(\ILAB0606.ILE0304.net2656 ));
  xci2_and3 _176__1 ( .a(\ILAB0606.net20227 ), .b(\ILAB0606.net22928 ), .c(\ILAB0606.net26797 ), .y(\ILAB0606.ILE0304.net0541 ));
  xci2_and3fft _177_ ( .a(\ILAB0606.net15799 ), .b(\ILAB0606.net16132 ), .c(\ILAB0606.net23357 ), .y(\ILAB0606.ILE0305.net2656 ));
  xci2_xnor2ft _178_ ( .a(\ILAB0606.net15548 ), .b(\ILAB0606.ILE0405.net01342 ), .y(\ILAB0606.ILE0405.net0541 ));
  xci2_and3 _179_ ( .a(\ILAB0606.ILE0107.net01342 ), .b(\ILAB0606.net17528 ), .c(\ILAB0606.ILE0506.net01339 ), .y(\ILAB0606.ILE0506.net2656 ));
  xci2_aoi21 _180_ ( .a(\ILAB0606.net20182 ), .b(\ILAB0606.net16114 ), .c(\ILAB0606.net26212 ), .y(\ILAB0606.ILE0404.net2656 ));
  xci2_and3 _181_ ( .a(\net14051<3> ), .b(\ILAB0606.net26214 ), .c(\ILAB0606.ILE0403.net01339 ), .y(\ILAB0606.ILE0403.net2656 ));
  xci2_and3 _181__1 ( .a(\net14051<3> ), .b(\ILAB0606.net26214 ), .c(\ILAB0606.ILE0403.net01339 ), .y(\ILAB0606.ILE0403.net0541 ));
  xci2_and3fft _182_ ( .a(\ILAB0606.net26213 ), .b(\ILAB0606.ILE0502.net01339 ), .c(\ILAB0606.net26464 ), .y(\ILAB0606.ILE0502.net2656 ));
  xci2_xnor2ft _183_ ( .a(\ILAB0606.net26258 ), .b(\ILAB0606.net17687 ), .y(\ILAB0606.ILE0503.net2656 ));
  xci2_and3 _184_ ( .a(\ILAB0606.ILE0107.net01342 ), .b(\ILAB0606.net17685 ), .c(\ILAB0606.net20137 ), .y(\ILAB0606.ILE0505.net2656 ));
  xci2_and3 _185_ ( .a(\net14047<6> ), .b(\net14047<3> ), .c(\ILAB0606.net20723 ), .y(\ILAB0606.ILE0501.net2656 ));
  xci2_and3 _185__1 ( .a(\net14047<6> ), .b(\net14047<3> ), .c(\ILAB0606.net20723 ), .y(\ILAB0606.ILE0501.net0541 ));
  xci2_aoi21 _186_ ( .a(\net14047<6> ), .b(\net14051<6> ), .c(\net14047<3> ), .y(\ILAB0606.ILE0401.net0541 ));
  xci2_and3fft _187_ ( .a(\net14047<1> ), .b(\ILAB0605.ILE0516.net01339 ), .c(\ILAB0605.ILE0516.net01342 ), .y(\ILAB0605.ILE0516.net2656 ));
  xci2_oai21 _188_ ( .a(\net14043<1> ), .b(\net14047<2> ), .c(\ILAB0605.net22099 ), .y(\ILAB0605.ILE0615.net2656 ));
  xci2_aoi21 _189_ ( .a(\net14043<2> ), .b(\ILAB0605.ILE0616.net01342 ), .c(\ILAB0605.net23964 ), .y(\ILAB0605.ILE0616.net2656 ));
  xci2_and3 _190_ ( .a(\net14043<0> ), .b(\ILAB0605.net24097 ), .c(\net14047<1> ), .y(\ILAB0605.ILE0614.net2656 ));
  xci2_and3 _190__1 ( .a(\net14043<0> ), .b(\ILAB0605.net24097 ), .c(\net14047<1> ), .y(\ILAB0605.ILE0614.net0541 ));
  xci2_aoi21 _191_ ( .a(\net14043<0> ), .b(\net14047<0> ), .c(\ILAB0605.ILE0514.net0558 ), .y(\ILAB0605.ILE0514.net2656 ));
  xci2_and3fft _192_ ( .a(\ILAB0605.ILE0513.net0562 ), .b(\ILAB0605.net23917 ), .c(\ILAB0605.net19354 ), .y(\ILAB0605.ILE0513.net2656 ));
  xci2_oai21 _193_ ( .a(\ILAB0605.ILE0411.net0562 ), .b(\ILAB0605.net22144 ), .c(\ILAB0605.net19892 ), .y(\ILAB0605.ILE0411.net2656 ));
  xci2_aoi21 _194_ ( .a(\ILAB0605.net23942 ), .b(\ILAB0605.net18112 ), .c(\ILAB0605.net16672 ), .y(\ILAB0605.ILE0410.net2656 ));
  xci2_ao21 _195_ ( .a(\ILAB0605.ILE0611.net01345 ), .b(\ILAB0605.net17077 ), .c(\ILAB0605.net18499 ), .y(\ILAB0605.ILE0611.net2656 ));
  xci2_nand2 _196_ ( .a(\ILAB0605.net20364 ), .b(\ILAB0605.ILE0513.net0562 ), .y(\ILAB0605.ILE0512.net2656 ));
  xci2_and3 _197_ ( .a(\ILAB0605.net16339 ), .b(\ILAB0605.net21444 ), .c(\ILAB0605.net18949 ), .y(\ILAB0605.ILE0612.net0541 ));
  xci2_aoi21 _198_ ( .a(\ILAB0605.ILE0412.net0562 ), .b(\ILAB0605.net22144 ), .c(\ILAB0605.ILE0412.net01339 ), .y(\ILAB0605.ILE0412.net2656 ));
  xci2_and3 _199_ ( .a(\ILAB0605.net19984 ), .b(\ILAB0605.net21467 ), .c(\ILAB0605.net22144 ), .y(\ILAB0605.ILE0413.net2656 ));
  xci2_and3 _199__1 ( .a(\ILAB0605.net19984 ), .b(\ILAB0605.net21467 ), .c(\ILAB0605.net22144 ), .y(\ILAB0605.ILE0413.net0541 ));
  xci2_and3fft _200_ ( .a(\net14018<6> ), .b(\ILAB0605.ILE0312.net0558 ), .c(\net14018<3> ), .y(\ILAB0605.ILE0312.net2656 ));
  xci2_oai21 _201_ ( .a(\ILAB0605.ILE0211.net0562 ), .b(\net14014<6> ), .c(\net14022<3> ), .y(\ILAB0605.ILE0211.net2656 ));
  xci2_aoi21 _202_ ( .a(\ILAB0605.net25899 ), .b(\net14014<6> ), .c(\ILAB0605.net21469 ), .y(\ILAB0605.ILE0311.net2656 ));
  xci2_aoi21 _203_ ( .a(\ILAB0605.net22299 ), .b(\net14014<6> ), .c(\ILAB0605.net23085 ), .y(\ILAB0605.ILE0213.net0541 ));
  xci2_and3 _204_ ( .a(\ILAB0605.net23897 ), .b(\ILAB0605.ILE0212.net01342 ), .c(\net14014<6> ), .y(\ILAB0605.ILE0212.net2656 ));
  xci2_and3 _204__1 ( .a(\ILAB0605.net23897 ), .b(\ILAB0605.ILE0212.net01342 ), .c(\net14014<6> ), .y(\ILAB0605.ILE0212.net0541 ));
  xci2_and3fft _205_ ( .a(\ILAB0605.ILE0112.net0562 ), .b(\net14018<1> ), .c(\net14018<4> ), .y(\ILAB0605.ILE0112.net2656 ));
  xci2_oai21 _206_ ( .a(\ILAB0605.ILE0111.net01345 ), .b(\ILAB0605.ILE0111.net0560 ), .c(\net14022<3> ), .y(\ILAB0605.ILE0111.net2656 ));
  xci2_aoi21 _207_ ( .a(\net14026<6> ), .b(\net14018<1> ), .c(\ILAB0605.net16807 ), .y(\ILAB0605.ILE0110.net2656 ));
  xci2_aoi21 _208_ ( .a(\ILAB0505.net24367 ), .b(\net14018<1> ), .c(\ILAB0505.ILE1612.net01339 ), .y(\ILAB0505.ILE1612.net2656 ));
  xci2_and3 _209_ ( .a(\ILAB0505.net22005 ), .b(\ILAB0505.net24367 ), .c(\net14018<1> ), .y(\ILAB0505.ILE1611.net2656 ));
  xci2_and3 _209__1 ( .a(\ILAB0505.net22005 ), .b(\ILAB0505.net24367 ), .c(\net14018<1> ), .y(\ILAB0505.ILE1611.net0541 ));
  xci2_and3fft _210_ ( .a(\net13659<3> ), .b(\ILAB0505.Clk_LAB<3> ), .c(\net13709<0> ), .y(\ILAB0505.ILE1512.net2656 ));
  xci2_oai21 _211_ ( .a(\ILAB0505.ILE1411.net01345 ), .b(\net13659<2> ), .c(\ILAB0505.net18067 ), .y(\ILAB0505.ILE1411.net2656 ));
  xci2_aoi21 _212_ ( .a(\net14018<0> ), .b(\ILAB0505.Clk_LAB<3> ), .c(\ILAB0505.net20409 ), .y(\ILAB0505.ILE1412.net2656 ));
  xci2_aoi21 _213_ ( .a(\ILAB0505.ILE1413.net01345 ), .b(\ILAB0505.Clk_LAB<3> ), .c(\ILAB0505.ILE1413.net01339 ), .y(\ILAB0505.ILE1413.net2656 ));
  xci2_and3 _214_ ( .a(\ILAB0505.net20115 ), .b(\ILAB0505.net22052 ), .c(\ILAB0505.Clk_LAB<3> ), .y(\ILAB0505.ILE1513.net2656 ));
  xci2_and3fft _215_ ( .a(\ILAB0505.net18364 ), .b(\ILAB0505.net19219 ), .c(\ILAB0505.net24682 ), .y(\ILAB0505.ILE1313.net2656 ));
  xci2_oa21 _216_ ( .a(\ILAB0505.net22050 ), .b(\net13713<5> ), .c(\net13709<0> ), .y(\ILAB0505.ILE1416.net2656 ));
  xci2_and2 _217_ ( .a(\net13717<4> ), .b(\ILAB0505.net19217 ), .y(\ILAB0505.ILE1316.net2656 ));
  xci2_and2 _217__1 ( .a(\net13717<4> ), .b(\ILAB0505.net19217 ), .y(\ILAB0505.ILE1316.net0541 ));
  xci2_and2ft _218_ ( .a(\ILAB0505.net20972 ), .b(\ILAB0505.net17914 ), .y(\ILAB0505.ILE1216.net2656 ));
  xci2_oai21 _219_ ( .a(\ILAB0505.net24302 ), .b(\ILAB0505.net23243 ), .c(\ILAB0506.net25067 ), .y(\ILAB0505.ILE1315.net2656 ));
  xci2_aoi21 _220_ ( .a(\ILAB0505.net24435 ), .b(\ILAB0505.ILE1215.net0560 ), .c(\ILAB0505.net24304 ), .y(\ILAB0505.ILE1215.net2656 ));
  xci2_ao21 _221_ ( .a(\ILAB0506.net16584 ), .b(\ILAB0506.ILE1201.net0560 ), .c(\ILAB0506.net15521 ), .y(\ILAB0506.ILE1201.net0541 ));
  xci2_and3 _222_ ( .a(\ILAB0505.net22050 ), .b(\net15119<0> ), .c(\net13705<0> ), .y(\ILAB0506.ILE1501.net2656 ));
  xci2_nand3 _223_ ( .a(\ILAB0505.net22050 ), .b(\net15119<0> ), .c(\net13705<0> ), .y(\ILAB0506.ILE1401.net2656 ));
  xci2_nand3 _223__1 ( .a(\ILAB0505.net22050 ), .b(\net15119<0> ), .c(\net13705<0> ), .y(\ILAB0506.ILE1401.net0541 ));
  xci2_and3 _224_ ( .a(\ILAB0506.net25067 ), .b(\ILAB0506.ILE1302.net01342 ), .c(\ILAB0506.ILE1302.net0558 ), .y(\ILAB0506.ILE1302.net2656 ));
  xci2_aoi21ttf _225_ ( .a(\ILAB0506.net26303 ), .b(\ILAB0506.net20857 ), .c(\ILAB0506.net20812 ), .y(\ILAB0506.ILE1403.net2656 ));
  xci2_aoi21ftf _226_ ( .a(\net13709<6> ), .b(\ILAB0506.net20814 ), .c(\net13709<3> ), .y(\ILAB0506.ILE1402.net2656 ));
  xci2_aoi21 _227_ ( .a(\ILAB0506.net25382 ), .b(\ILAB0506.net20857 ), .c(\ILAB0506.net25384 ), .y(\ILAB0506.ILE1504.net0541 ));
  xci2_and3 _228_ ( .a(\ILAB0506.ILE1503.net01345 ), .b(\ILAB0506.ILE1503.net0560 ), .c(\ILAB0506.net20857 ), .y(\ILAB0506.ILE1503.net2656 ));
  xci2_and3fft _229_ ( .a(\ILAB0506.ILE1603.net01345 ), .b(\ILAB0506.net15484 ), .c(\net15111<3> ), .y(\ILAB0506.ILE1603.net2656 ));
  xci2_oai21 _230_ ( .a(\ILAB0505.net24257 ), .b(\net13705<3> ), .c(\ILAB0506.net20812 ), .y(\ILAB0505.ILE1615.net2656 ));
  xci2_aoi21 _231_ ( .a(\ILAB0505.net22815 ), .b(\ILAB0505.net19642 ), .c(\net13659<6> ), .y(\ILAB0505.ILE1515.net2656 ));
  xci2_ao21 _232_ ( .a(\ILAB0505.ILE1516.net01345 ), .b(\net13705<3> ), .c(\net13705<1> ), .y(\ILAB0505.ILE1516.net0541 ));
  xci2_nand3 _233_ ( .a(\ILAB0505.net24257 ), .b(\net13705<5> ), .c(\net13705<6> ), .y(\ILAB0505.ILE1616.net2656 ));
  xci2_and3 _234_ ( .a(\ILAB0506.net20812 ), .b(\ILAB0506.ILE1601.net01342 ), .c(\net13701<5> ), .y(\ILAB0506.ILE1601.net0541 ));
  xci2_xnor2 _235_ ( .a(\ILAB0605.ILE0116.net0558 ), .b(\net14002<0> ), .y(\ILAB0605.ILE0116.net2656 ));
  xci2_and2 _236_ ( .a(\net15111<3> ), .b(\ILAB0605.net21892 ), .y(\ILAB0605.ILE0115.net2656 ));
  xci2_aoi21ftf _237_ ( .a(\ILAB0506.net24952 ), .b(\ILAB0506.net18049 ), .c(\ILAB0506.Clk_LAB<3> ), .y(\ILAB0506.ILE1112.net2656 ));
  xci2_or2ft _238_ ( .a(\ILAB0506.net23537 ), .b(\ILAB0506.net22657 ), .y(\ILAB0506.ILE1014.net2656 ));
  xci2_or2ft _238__1 ( .a(\ILAB0506.net23537 ), .b(\ILAB0506.net22657 ), .y(\ILAB0506.ILE1014.net0541 ));
  xci2_and2 _239_ ( .a(\ILAB0506.net21759 ), .b(\ILAB0506.ILE1113.net01339 ), .y(\ILAB0506.ILE1113.net2656 ));
  xci2_aoi21ftf _240_ ( .a(\ILAB0506.ILE1013.net01345 ), .b(\ILAB0506.net24862 ), .c(\ILAB0506.Clk_LAB<3> ), .y(\ILAB0506.ILE1013.net2656 ));
  xci2_and3 _241_ ( .a(\ILAB0506.net24952 ), .b(\ILAB0506.net21690 ), .c(\ILAB0506.net24682 ), .y(\ILAB0506.ILE1012.net2656 ));
  xci2_and3 _241__1 ( .a(\ILAB0506.net24952 ), .b(\ILAB0506.net21690 ), .c(\ILAB0506.net24682 ), .y(\ILAB0506.ILE1012.net0541 ));
  xci2_nand2 _242_ ( .a(\ILAB0506.net23537 ), .b(\ILAB0506.net18922 ), .y(\ILAB0506.ILE0915.net2656 ));
  xci2_and2ft _243_ ( .a(\ILAB0506.ILE0913.net0562 ), .b(\ILAB0506.net21424 ), .y(\ILAB0506.ILE0913.net2656 ));
  xci2_or2 _244_ ( .a(\ILAB0506.ILE0813.net01345 ), .b(\ILAB0506.net21692 ), .y(\ILAB0506.ILE0813.net2656 ));
  xci2_or3ftt _245_ ( .a(\ILAB0506.net23539 ), .b(\ILAB0506.net18967 ), .c(\ILAB0506.net25493 ), .y(\ILAB0506.ILE0914.net2656 ));
  xci2_and3 _246_ ( .a(\ILAB0506.ILE0716.net01345 ), .b(\ILAB0506.net22549 ), .c(\ILAB0506.net23494 ), .y(\ILAB0506.ILE0713.net2656 ));
  xci2_aoi21ftf _247_ ( .a(\ILAB0506.ILE0712.net01345 ), .b(\ILAB0506.net23494 ), .c(\ILAB0506.Clk_LAB<3> ), .y(\ILAB0506.ILE0712.net2656 ));
  xci2_nand3 _248_ ( .a(\ILAB0506.ILE0613.net0562 ), .b(\ILAB0506.net19687 ), .c(\ILAB0506.net21694 ), .y(\ILAB0506.ILE0613.net2656 ));
  xci2_and2 _249_ ( .a(\ILAB0506.net19939 ), .b(\ILAB0506.net21443 ), .y(\ILAB0506.ILE0612.net2656 ));
  xci2_aoi21ftf _250_ ( .a(\ILAB0506.net20389 ), .b(\ILAB0506.net19354 ), .c(\ILAB0506.Clk_LAB<3> ), .y(\ILAB0506.ILE0311.net2656 ));
  xci2_or2ft _251_ ( .a(\ILAB0506.net20387 ), .b(\ILAB0506.net19354 ), .y(\ILAB0506.ILE0312.net2656 ));
  xci2_or2ft _251__1 ( .a(\ILAB0506.net20387 ), .b(\ILAB0506.net19354 ), .y(\ILAB0506.ILE0312.net0541 ));
  xci2_and2 _252_ ( .a(\ILAB0506.net21514 ), .b(\ILAB0506.ILE0411.net01339 ), .y(\ILAB0506.ILE0411.net2656 ));
  xci2_aoi21ftf _253_ ( .a(\ILAB0506.net19084 ), .b(\net14773<6> ), .c(\ILAB0506.Clk_LAB<3> ), .y(\ILAB0506.ILE0412.net2656 ));
  xci2_or3fft _254_ ( .a(\ILAB0506.net20387 ), .b(\ILAB0506.net19082 ), .c(\ILAB0506.net19354 ), .y(\ILAB0506.ILE0313.net2656 ));
  xci2_and2 _255_ ( .a(\ILAB0506.net19014 ), .b(\ILAB0506.net19984 ), .y(\ILAB0506.ILE0413.net0541 ));
  xci2_aoi21ftf _256_ ( .a(\ILAB0506.net19804 ), .b(\net14810<0> ), .c(\ILAB0506.Clk_LAB<3> ), .y(\ILAB0506.ILE0314.net2656 ));
  xci2_nor2ft _257_ ( .a(\ILAB0506.ILE0415.net0562 ), .b(\ILAB0506.net24819 ), .y(\ILAB0506.ILE0415.net2656 ));
  xci2_and2ft _258_ ( .a(\ILAB0506.net26078 ), .b(\ILAB0506.net22414 ), .y(\ILAB0506.ILE0414.net2656 ));
  xci2_xnor2 _259_ ( .a(\ILAB0506.ILE0515.net0558 ), .b(\ILAB0506.net22099 ), .y(\ILAB0506.ILE0515.net2656 ));
  xci2_and2ft _260_ ( .a(\ILAB0506.net22189 ), .b(\ILAB0506.Clk_LAB<3> ), .y(\ILAB0506.ILE0615.net2656 ));
  xci2_xnor2 _261_ ( .a(\ILAB0606.net16249 ), .b(\ILAB0606.net16294 ), .y(\ILAB0606.ILE1209.net2656 ));
  xci2_and2 _262_ ( .a(\ILAB0606.ILE1016.net01339 ), .b(\ILAB0606.net16292 ), .y(\ILAB0606.ILE1109.net2656 ));
  xci2_nand3fft _263_ ( .a(\ILAB0606.net16222 ), .b(\ILAB0606.net24682 ), .c(\ILAB0606.net24728 ), .y(\ILAB0606.ILE1312.net2656 ));
  xci2_nand3fft _263__1 ( .a(\ILAB0606.net16222 ), .b(\ILAB0606.net24682 ), .c(\ILAB0606.net24728 ), .y(\ILAB0606.ILE1312.net0541 ));
  xci2_oa21ftt _264_ ( .a(\ILAB0606.net21758 ), .b(\ILAB0606.net21242 ), .c(\ILAB0606.net24728 ), .y(\ILAB0606.ILE1212.net0541 ));
  xci2_xnor2ft _265_ ( .a(\ILAB0606.ILE1410.net01339 ), .b(\ILAB0606.net24032 ), .y(\ILAB0606.ILE1410.net2656 ));
  xci2_mux2h _266_ ( .a(\ILAB0606.ILE1111.net0562 ), .b(\ILAB0606.net24034 ), .s(\ILAB0606.net23040 ), .y(\ILAB0606.ILE1111.net2656 ));
  xci2_and2 _267_ ( .a(\ILAB0606.ILE1016.net01339 ), .b(\ILAB0606.net16358 ), .y(\ILAB0606.ILE1110.net2656 ));
  xci2_or3fft _268_ ( .a(\ILAB0606.net18092 ), .b(\ILAB0606.net24729 ), .c(\ILAB0606.net15349 ), .y(\ILAB0606.ILE1211.net2656 ));
  xci2_and3 _269_ ( .a(\net14936<1> ), .b(\ILAB0606.net24075 ), .c(\ILAB0606.ILE1411.net01339 ), .y(\ILAB0606.ILE1412.net2656 ));
  xci2_aoi21ftf _270_ ( .a(\ILAB0606.net21784 ), .b(\ILAB0606.net19399 ), .c(\ILAB0606.ILE1016.net01339 ), .y(\ILAB0606.ILE1112.net2656 ));
  xci2_aoi21ftf _271_ ( .a(\ILAB0606.net24684 ), .b(\net15018<2> ), .c(\ILAB0606.net23018 ), .y(\ILAB0606.ILE1311.net2656 ));
  xci2_and3 _272_ ( .a(\ILAB0606.ILE1213.net01345 ), .b(\ILAB0606.net22567 ), .c(\ILAB0606.ILE1213.net0558 ), .y(\ILAB0606.ILE1213.net2656 ));
  xci2_nand2ft _273_ ( .a(\ILAB0606.net23017 ), .b(\ILAB0606.ILE1411.net01339 ), .y(\ILAB0606.ILE1411.net2656 ));
  xci2_nand2ft _274_ ( .a(\net14916<4> ), .b(\net15068<2> ), .y(\ILAB0606.ILE1615.net2656 ));
  xci2_nand2ft _274__1 ( .a(\net14916<4> ), .b(\net15068<2> ), .y(\ILAB0606.ILE1615.net0541 ));
  xci2_xnor2ft _275_ ( .a(\ILAB0606.net22054 ), .b(\ILAB0606.net19397 ), .y(\ILAB0606.ILE1214.net2656 ));
  xci2_nand2ft _276_ ( .a(\ILAB0606.net23539 ), .b(\ILAB0606.net23449 ), .y(\ILAB0606.ILE1014.net2656 ));
  xci2_aoi21ftf _277_ ( .a(\ILAB0606.net21109 ), .b(\ILAB0606.net24862 ), .c(\ILAB0606.ILE1016.net01339 ), .y(\ILAB0606.ILE1013.net0541 ));
  xci2_or2 _278_ ( .a(\ILAB0606.net24075 ), .b(\ILAB0606.net20993 ), .y(\ILAB0606.ILE1413.net2656 ));
  xci2_ao21ftt _279_ ( .a(\ILAB0606.net19372 ), .b(\net15068<0> ), .c(\ILAB0606.net22772 ), .y(\ILAB0606.ILE1415.net0541 ));
  xci2_ao21ttf _280_ ( .a(\ILAB0606.net16020 ), .b(\ILAB0606.net18338 ), .c(\ILAB0606.net20993 ), .y(\ILAB0606.ILE1513.net2656 ));
  xci2_oai21ttf _281_ ( .a(\ILAB0606.net19373 ), .b(\ILAB0606.net24075 ), .c(\ILAB0606.net22054 ), .y(\ILAB0606.ILE1414.net2656 ));
  xci2_oai21ttf _281__1 ( .a(\ILAB0606.net19373 ), .b(\ILAB0606.net24075 ), .c(\ILAB0606.net22054 ), .y(\ILAB0606.ILE1414.net0541 ));
  xci2_mux2h _282_ ( .a(\ILAB0606.net24390 ), .b(\net14928<1> ), .s(\net14928<0> ), .y(\ILAB0606.ILE1511.net2656 ));
  xci2_ao21ftt _283_ ( .a(\ILAB0606.net22054 ), .b(\ILAB0606.net19643 ), .c(\ILAB0606.net21262 ), .y(\ILAB0606.ILE1514.net2656 ));
  xci2_oai21 _284_ ( .a(\ILAB0606.net18338 ), .b(\ILAB0606.net20993 ), .c(\ILAB0606.net21083 ), .y(\ILAB0606.ILE1613.net2656 ));
  xci2_oai21 _284__1 ( .a(\ILAB0606.net18338 ), .b(\ILAB0606.net20993 ), .c(\ILAB0606.net21083 ), .y(\ILAB0606.ILE1613.net0541 ));
  xci2_nand2ft _285_ ( .a(\ILAB0606.ILE1515.net01345 ), .b(\net15064<0> ), .y(\ILAB0606.ILE1515.net0541 ));
  xci2_ao21ftt _286_ ( .a(\ILAB0606.net21354 ), .b(\ILAB0606.net24390 ), .c(\ILAB0606.net21218 ), .y(\ILAB0606.ILE1512.net2656 ));
  xci2_nand2 _287_ ( .a(\net14920<6> ), .b(\ILAB0706.net22320 ), .y(\ILAB0706.ILE0113.net0541 ));
  xci2_xnor2ft _288_ ( .a(\ILAB0606.net21354 ), .b(\net14932<5> ), .y(\ILAB0606.ILE1612.net2656 ));
  xci2_aoi21ftf _289_ ( .a(\net14916<1> ), .b(\ILAB0606.net20092 ), .c(\net14916<3> ), .y(\ILAB0606.ILE1614.net2656 ));
  xci2_aoi21ftf _289__1 ( .a(\net14916<1> ), .b(\ILAB0606.net20092 ), .c(\net14916<3> ), .y(\ILAB0606.ILE1614.net0541 ));
  xci2_nand2 _290_ ( .a(\ILAB0706.Clk_LAB<0> ), .b(\net14916<6> ), .y(\ILAB0706.ILE0114.net0541 ));
  xci2_or2 _291_ ( .a(\ILAB0606.net21011 ), .b(\ILAB0606.net21219 ), .y(\ILAB0606.ILE1313.net2656 ));
  xci2_or2ft _292_ ( .a(\net14932<4> ), .b(\net14928<1> ), .y(\ILAB0606.ILE1611.net0541 ));
  xci2_nand2 _293_ ( .a(\net14912<6> ), .b(\ILAB0706.Clk_LAB<1> ), .y(\ILAB0706.ILE0115.net0541 ));
  xci2_dff _294_ ( .d(\net15022<6> ), .clk(\ILAB0606.net18589 ), .q(\ILAB0606.ILE0207.net2656 ));
  xci2_dff _295_ ( .d(\net15099<4> ), .clk(\ILAB0606.ILE0106.net01342 ), .q(\ILAB0606.ILE0106.net2656 ));
  xci2_dff _295__1 ( .d(\net15099<4> ), .clk(\ILAB0606.ILE0106.net01342 ), .q(\ILAB0606.ILE0106.net0541 ));
  xci2_dff _296_ ( .d(\ILAB0606.net23334 ), .clk(\ILAB0606.net17552 ), .q(\ILAB0606.ILE0306.net2656 ));
  xci2_dff _296__1 ( .d(\ILAB0606.net23334 ), .clk(\ILAB0606.net17552 ), .q(\ILAB0606.ILE0306.net0541 ));
  xci2_dff _297_ ( .d(\net15022<5> ), .clk(\ILAB0606.net18589 ), .q(\ILAB0606.ILE0406.net2656 ));
  xci2_dff _298_ ( .d(\net15022<1> ), .clk(\ILAB0506.ILE1604.net0560 ), .q(\ILAB0606.ILE0402.net2656 ));
  xci2_dff _298__1 ( .d(\net15022<1> ), .clk(\ILAB0506.ILE1604.net0560 ), .q(\ILAB0606.ILE0402.net0541 ));
  xci2_dff _299_ ( .d(\ILAB0606.net20632 ), .clk(\ILAB0606.Clk_LAB<2> ), .q(\ILAB0606.ILE0504.net2656 ));
  xci2_dff _300_ ( .d(\ILAB0605.net19057 ), .clk(\ILAB0605.net20362 ), .q(\ILAB0605.ILE0515.net2656 ));
  xci2_dff _300__1 ( .d(\ILAB0605.net19057 ), .clk(\ILAB0605.net20362 ), .q(\ILAB0605.ILE0515.net0541 ));
  xci2_dff _301_ ( .d(\net14043<4> ), .clk(\ILAB0606.ILE0601.net01342 ), .q(\ILAB0606.ILE0601.net2656 ));
  xci2_dff _302_ ( .d(\ILAB0605.net25519 ), .clk(\ILAB0605.Clk_LAB<2> ), .q(\ILAB0605.ILE0613.net2656 ));
  xci2_dff _302__1 ( .d(\ILAB0605.net25519 ), .clk(\ILAB0605.Clk_LAB<2> ), .q(\ILAB0605.ILE0613.net0541 ));
  xci2_dff _303_ ( .d(\ILAB0605.net23629 ), .clk(\ILAB0605.ILE0113.net01342 ), .q(\ILAB0605.ILE0510.net2656 ));
  xci2_dff _303__1 ( .d(\ILAB0605.net23629 ), .clk(\ILAB0605.ILE0113.net01342 ), .q(\ILAB0605.ILE0510.net0541 ));
  xci2_dff _304_ ( .d(\ILAB0605.ILE0711.net01345 ), .clk(\ILAB0605.net18319 ), .q(\ILAB0605.ILE0711.net2656 ));
  xci2_dff _305_ ( .d(\ILAB0605.net24909 ), .clk(\ILAB0605.net18319 ), .q(\ILAB0605.ILE0313.net2656 ));
  xci2_dff _305__1 ( .d(\ILAB0605.net24909 ), .clk(\ILAB0605.net18319 ), .q(\ILAB0605.ILE0313.net0541 ));
  xci2_dff _306_ ( .d(\ILAB0605.net25852 ), .clk(\ILAB0605.ILE0113.net01342 ), .q(\ILAB0605.ILE0310.net2656 ));
  xci2_dff _306__1 ( .d(\ILAB0605.net25852 ), .clk(\ILAB0605.ILE0113.net01342 ), .q(\ILAB0605.ILE0310.net0541 ));
  xci2_dff _307_ ( .d(\ILAB0605.net21894 ), .clk(\ILAB0605.ILE0113.net01342 ), .q(\ILAB0605.ILE0113.net2656 ));
  xci2_dff _307__1 ( .d(\ILAB0605.net21894 ), .clk(\ILAB0605.ILE0113.net01342 ), .q(\ILAB0605.ILE0113.net0541 ));
  xci2_dff _308_ ( .d(\net14026<0> ), .clk(\ILAB0505.ILE1610.net0560 ), .q(\ILAB0505.ILE1610.net2656 ));
  xci2_dff _308__1 ( .d(\net14026<0> ), .clk(\ILAB0505.ILE1610.net0560 ), .q(\ILAB0505.ILE1610.net0541 ));
  xci2_dff _309_ ( .d(\ILAB0505.net19552 ), .clk(\net14026<2> ), .q(\ILAB0505.ILE1511.net2656 ));
  xci2_dff _309__1 ( .d(\ILAB0505.net19552 ), .clk(\net14026<2> ), .q(\ILAB0505.ILE1511.net0541 ));
  xci2_dff _310_ ( .d(\ILAB0505.net19399 ), .clk(\ILAB0505.net21847 ), .q(\ILAB0505.ILE1312.net2656 ));
  xci2_dff _310__1 ( .d(\ILAB0505.net19399 ), .clk(\ILAB0505.net21847 ), .q(\ILAB0505.ILE1312.net0541 ));
  xci2_dff _311_ ( .d(\ILAB0505.net20994 ), .clk(\ILAB0605.ILE0113.net01342 ), .q(\ILAB0505.ILE1314.net2656 ));
  xci2_dff _311__1 ( .d(\ILAB0505.net20994 ), .clk(\ILAB0605.ILE0113.net01342 ), .q(\ILAB0505.ILE1314.net0541 ));
  xci2_dff _312_ ( .d(\ILAB0505.net21352 ), .clk(\ILAB0505.ILE1610.net0560 ), .q(\ILAB0505.ILE1214.net2656 ));
  xci2_dff _313_ ( .d(\ILAB0505.net24439 ), .clk(\ILAB0506.ILE1101.net01339 ), .q(\ILAB0505.ILE1115.net2656 ));
  xci2_dff _314_ ( .d(\ILAB0506.net26554 ), .clk(\net13717<1> ), .q(\ILAB0506.ILE1202.net0541 ));
  xci2_dff _315_ ( .d(\ILAB0506.net26302 ), .clk(\ILAB0506.ILE1604.net0560 ), .q(\ILAB0506.ILE1404.net2656 ));
  xci2_dff _315__1 ( .d(\ILAB0506.net26302 ), .clk(\ILAB0506.ILE1604.net0560 ), .q(\ILAB0506.ILE1404.net0541 ));
  xci2_dff _316_ ( .d(\ILAB0506.net15459 ), .clk(\ILAB0506.ILE1604.net0560 ), .q(\ILAB0506.ILE1604.net2656 ));
  xci2_dff _316__1 ( .d(\ILAB0506.net15459 ), .clk(\ILAB0506.ILE1604.net0560 ), .q(\ILAB0506.ILE1604.net0541 ));
  xci2_dff _317_ ( .d(\ILAB0505.net22819 ), .clk(\ILAB0605.ILE0115.net01342 ), .q(\ILAB0505.ILE1415.net2656 ));
  xci2_dff _317__1 ( .d(\ILAB0505.net22819 ), .clk(\ILAB0605.ILE0115.net01342 ), .q(\ILAB0505.ILE1415.net0541 ));
  xci2_dff _318_ ( .d(\ILAB0506.Clk_LAB<1> ), .clk(\ILAB0506.Clk_LAB<2> ), .q(\ILAB0506.ILE1502.net2656 ));
  xci2_dff _319_ ( .d(\ILAB0605.net24615 ), .clk(\net14006<5> ), .q(\ILAB0605.ILE0215.net2656 ));
  xci2_dff _319__1 ( .d(\ILAB0605.net24615 ), .clk(\net14006<5> ), .q(\ILAB0605.ILE0215.net0541 ));
  xci2_dff _320_ ( .d(\ILAB0506.net21534 ), .clk(\ILAB0507.ILE1101.net01339 ), .q(\ILAB0506.ILE1114.net2656 ));
  xci2_dff _321_ ( .d(\ILAB0506.net25312 ), .clk(\ILAB0506.Clk_LAB<2> ), .q(\ILAB0506.ILE0912.net2656 ));
  xci2_dff _321__1 ( .d(\ILAB0506.net25312 ), .clk(\ILAB0506.Clk_LAB<2> ), .q(\ILAB0506.ILE0912.net0541 ));
  xci2_dff _322_ ( .d(\ILAB0506.net19959 ), .clk(\ILAB0507.ILE0701.net01339 ), .q(\ILAB0506.ILE0714.net2656 ));
  xci2_dff _322__1 ( .d(\ILAB0506.net19959 ), .clk(\ILAB0507.ILE0701.net01339 ), .q(\ILAB0506.ILE0714.net0541 ));
  xci2_dff _323_ ( .d(\ILAB0506.net24098 ), .clk(\ILAB0506.Clk_LAB<2> ), .q(\ILAB0506.ILE0611.net2656 ));
  xci2_dff _323__1 ( .d(\ILAB0506.net24098 ), .clk(\ILAB0506.Clk_LAB<2> ), .q(\ILAB0506.ILE0611.net0541 ));
  xci2_dff _324_ ( .d(\ILAB0506.net18499 ), .clk(\ILAB0506.Clk_LAB<2> ), .q(\ILAB0506.ILE0511.net2656 ));
  xci2_dff _325_ ( .d(\ILAB0506.ILE0512.net01345 ), .clk(\ILAB0506.Clk_LAB<2> ), .q(\ILAB0506.ILE0512.net2656 ));
  xci2_dff _326_ ( .d(\ILAB0506.net18904 ), .clk(\ILAB0507.ILE0501.net01339 ), .q(\ILAB0506.ILE0514.net2656 ));
  xci2_dff _326__1 ( .d(\ILAB0506.net18904 ), .clk(\ILAB0507.ILE0501.net01339 ), .q(\ILAB0506.ILE0514.net0541 ));
  xci2_dff _327_ ( .d(\ILAB0506.net21442 ), .clk(\ILAB0507.ILE0601.net01339 ), .q(\ILAB0506.ILE0614.net2656 ));
  xci2_dff _327__1 ( .d(\ILAB0506.net21442 ), .clk(\ILAB0507.ILE0601.net01339 ), .q(\ILAB0506.ILE0614.net0541 ));
  xci2_dff _328_ ( .d(\ILAB0606.net18049 ), .clk(\ILAB0606.ILE1609.net0562 ), .q(\ILAB0606.ILE1309.net2656 ));
  xci2_dff _328__1 ( .d(\ILAB0606.net18049 ), .clk(\ILAB0606.ILE1609.net0562 ), .q(\ILAB0606.ILE1309.net0541 ));
  xci2_dff _329_ ( .d(\ILAB0606.net24079 ), .clk(\ILAB0606.ILE1609.net0562 ), .q(\ILAB0606.ILE1210.net2656 ));
  xci2_dff _330_ ( .d(\ILAB0606.net17122 ), .clk(\ILAB0606.ILE1610.net0560 ), .q(\ILAB0606.ILE1310.net2656 ));
  xci2_dff _330__1 ( .d(\ILAB0606.net17122 ), .clk(\ILAB0606.ILE1610.net0560 ), .q(\ILAB0606.ILE1310.net0541 ));
  xci2_dff _331_ ( .d(\ILAB0606.ILE1114.net01345 ), .clk(\ILAB0607.ILE1101.net01339 ), .q(\ILAB0606.ILE1114.net2656 ));
  xci2_dff _331__1 ( .d(\ILAB0606.ILE1114.net01345 ), .clk(\ILAB0607.ILE1101.net01339 ), .q(\ILAB0606.ILE1114.net0541 ));
  mux2i_P_UCCLAB \IIO30.I7.I27  ( .d0(\IIO30.I7.net209 ), .d1(GND), .sl0(GND), .x(\IIO30.I7.net0151 ));
  mux2i_P_UCCLAB \IIO30.I7.I25  ( .d0(\IIO30.I7.net209 ), .d1(GND), .sl0(GND), .x(\IIO30.I7.net0153 ));
  invtd52_AVDD \IIO30.I7.I8  ( .a(\IIO30.I7.net0151 ), .en(VDD), .x(\LongBus_30<0> ));
  invtd52_AVDD \IIO30.I7.I26  ( .a(\IIO30.I7.net0153 ), .en(VDD), .x(\LongBus_31<8> ));
  buftd52C_UCCLAB \I1817.I62895  ( .a(\LongBus_30<0> ), .en(VDD), .x(\net8293<15> ));
  buftd52C_UCCLAB \I1818.I18  ( .a(\LongBus_31<8> ), .en(VDD), .x(\net8305<7> ));
  buftd52_UCCLAB \ILAB0604.I4772.I62895  ( .a(\net8293<15> ), .en(VDD), .x(\LongBus_10<0> ));
  buftd52_UCCLAB \ILAB0604.I4775.I62895  ( .a(\net8293<15> ), .en(VDD), .x(\LongBus_11<0> ));
  buftd52_UCCLAB \ILAB0504.I4801.I18  ( .a(\net8305<7> ), .en(VDD), .x(\LongBus_9<8> ));
  buftd52C_UCCLAB \I1839.I19  ( .a(\LongBus_9<8> ), .en(VDD), .x(\LongBus_50<8> ));
  buftd52C_UCCLAB \I1849.I1  ( .a(\LongBus_10<0> ), .en(VDD), .x(\LongBus_49<0> ));
  buftd52C_UCCLAB \I1848.I1  ( .a(\LongBus_11<0> ), .en(VDD), .x(\LongBus_48<0> ));
  buftd52_UCCLAB \ILAB0507.I4775.I19  ( .a(\LongBus_50<8> ), .en(VDD), .x(\net8308<7> ));
  buftd52_UCCLAB \ILAB0506.I4775.I19  ( .a(\LongBus_50<8> ), .en(VDD), .x(\net8314<7> ));
  inv_4_UCCLAB \ILAB0506.ILE1604.I711  ( .a(\LongBus_50<8> ), .x(\ILAB0506.ILE1604.net0560 ));
  inv_4_UCCLAB \ILAB0505.ILE1610.I711  ( .a(\LongBus_50<8> ), .x(\ILAB0505.ILE1610.net0560 ));
  inv_4_UCCLAB \ILAB0606.ILE0106.I713  ( .a(\LongBus_49<0> ), .x(\ILAB0606.ILE0106.net01342 ));
  inv_4_UCCLAB \ILAB0605.ILE0113.I713  ( .a(\LongBus_49<0> ), .x(\ILAB0605.ILE0113.net01342 ));
  inv_4_UCCLAB \ILAB0606.ILE0601.I713  ( .a(\net8314<7> ), .x(\ILAB0606.ILE0601.net01342 ));
  inv_4_UCCLAB \ILAB0606.ILE1609.I712  ( .a(\LongBus_48<0> ), .x(\ILAB0606.ILE1609.net0562 ));
  inv_4_UCCLAB \ILAB0607.ILE1101.I715  ( .a(\net8308<7> ), .x(\ILAB0607.ILE1101.net01339 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0106.Ivo2  ( .en(GND), .in(\ILAB0606.ILE0106.net01342 ), .out(\ILAB0606.net17552 ));
  buftd52_UCCLAB \ILAB0504.I4775.I62895  ( .a(\net8293<15> ), .en(VDD), .x(\LongBus_9<0> ));
  buftd52_UCCLAB \ILAB0604.I4773.I18  ( .a(\net8305<7> ), .en(VDD), .x(\LongBus_10<8> ));
  buftd52C_UCCLAB \I1839.I1  ( .a(\LongBus_9<0> ), .en(VDD), .x(\LongBus_50<0> ));
  buftd52C_UCCLAB \I1849.I19  ( .a(\LongBus_10<8> ), .en(VDD), .x(\LongBus_49<8> ));
  buftd52_UCCLAB \ILAB0507.I4775.I1  ( .a(\LongBus_50<0> ), .en(VDD), .x(\net8308<15> ));
  inv_4_UCCLAB \ILAB0506.ILE1605.I711  ( .a(\LongBus_50<0> ), .x(\ILAB0506.ILE1605.net0560 ));
  inv_4_UCCLAB \ILAB0606.ILE1610.I711  ( .a(\LongBus_48<0> ), .x(\ILAB0606.ILE1610.net0560 ));
  inv_4_UCCLAB \ILAB0506.ILE1101.I715  ( .a(\net8314<7> ), .x(\ILAB0506.ILE1101.net01339 ));
  inv_4_UCCLAB \ILAB0507.ILE0601.I715  ( .a(\net8308<15> ), .x(\ILAB0507.ILE0601.net01339 ));
  inv_4_UCCLAB \ILAB0507.ILE0701.I715  ( .a(\net8308<15> ), .x(\ILAB0507.ILE0701.net01339 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0113.Ivo1  ( .en(GND), .in(\ILAB0605.ILE0113.net01342 ), .out(\ILAB0605.net18319 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0206.Ivo1  ( .en(GND), .in(\ILAB0606.ILE0106.net01342 ), .out(\ILAB0606.net18589 ));
  inv_8_UCCLAB \ILAB0506.ILE1605.I666  ( .a(\ILAB0506.ILE1605.net0560 ), .x(\ILAB0506.net25376 ));
  buftd4_UCCLAB \ILAB0506.I222  ( .a(\ILAB0506.net25376 ), .en(VDD), .x(\ILAB0506.net27128 ));
  mux2p_2_UCCLAB \ILAB0506.I5605.I2  ( .d0(\ILAB0506.net27128 ), .d1(GND), .s0(GND), .x(\ILAB0506.I5605.net33 ));
  invd16_seth_UCCLAB \ILAB0506.I5605.I3  ( .a(\ILAB0506.I5605.net33 ), .c(VDD), .x(\ILAB0506.Clk_int<2> ));
  mux2d1i_1_P_UCCLAB \ILAB0506.I5366.I80  ( .d0(\ILAB0506.Clk_int<2> ), .d1i(GND), .sl0(GND), .x(\ILAB0506.I5366.net0106 ));
  invd52_UCCLAB \ILAB0506.I5366.I76  ( .a(\ILAB0506.I5366.net0106 ), .x(\ILAB0506.net15299<1> ));
  invd32_UCCLAB \ILAB0506.I5591.I1  ( .a(\ILAB0506.net15299<1> ), .x(\ILAB0506.Clk_LAB<2> ));
  buftd52_UCCLAB \ILAB0505.I4801.I1  ( .a(\LongBus_50<0> ), .en(VDD), .x(\net8290<15> ));
  inv_4_UCCLAB \ILAB0605.ILE0115.I713  ( .a(\LongBus_49<8> ), .x(\ILAB0605.ILE0115.net01342 ));
  inv_4_UCCLAB \ILAB0606.ILE1609.I710  ( .a(\LongBus_48<0> ), .x(\ILAB0606.ILE1609.net0558 ));
  inv_4_UCCLAB \ILAB0507.ILE1101.I715  ( .a(\net8308<15> ), .x(\ILAB0507.ILE1101.net01339 ));
  inv_4_UCCLAB \ILAB0507.ILE0501.I715  ( .a(\net8308<15> ), .x(\ILAB0507.ILE0501.net01339 ));
  inv_4_UCCLAB \ILAB0505.ILE1316.I713  ( .a(\net8290<15> ), .x(\ILAB0505.ILE1316.net01342 ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1510.Ivo2  ( .en(GND), .in(\ILAB0505.ILE1610.net0560 ), .out(\net14026<2> ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1214.Iho1  ( .en(GND), .in(\ILAB0505.ILE1610.net0560 ), .out(\net13717<1> ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1615.Ivo2  ( .en(GND), .in(\ILAB0605.ILE0115.net01342 ), .out(\net14006<5> ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1312.Ihi7  ( .en(GND), .in(\ILAB0505.ILE1316.net01342 ), .out(\ILAB0505.net21847 ));
  inv_8_UCCLAB \ILAB0606.ILE1609.I666  ( .a(\ILAB0606.ILE1609.net0558 ), .x(\ILAB0606.net21641 ));
  buftd4_UCCLAB \ILAB0606.I206  ( .a(\ILAB0606.net21641 ), .en(VDD), .x(\ILAB0606.net015238 ));
  mux2p_2_UCCLAB \ILAB0606.I5605.I2  ( .d0(GND), .d1(\ILAB0606.net015238 ), .s0(VDD), .x(\ILAB0606.I5605.net33 ));
  invd16_seth_UCCLAB \ILAB0606.I5605.I3  ( .a(\ILAB0606.I5605.net33 ), .c(VDD), .x(\ILAB0606.Clk_int<2> ));
  mux2d1i_1_P_UCCLAB \ILAB0606.I5366.I80  ( .d0(\ILAB0606.Clk_int<2> ), .d1i(GND), .sl0(GND), .x(\ILAB0606.I5366.net0106 ));
  invd52_UCCLAB \ILAB0606.I5366.I76  ( .a(\ILAB0606.I5366.net0106 ), .x(\ILAB0606.net15299<1> ));
  invd32_UCCLAB \ILAB0606.I5591.I1  ( .a(\ILAB0606.net15299<1> ), .x(\ILAB0606.Clk_LAB<2> ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0511.Iho1  ( .en(GND), .in(\ILAB0605.ILE0113.net01342 ), .out(\ILAB0605.net20362 ));
  inv_4_UCCLAB \ILAB1004.ILE1616.I713  ( .a(\LongBus_31<8> ), .x(\ILAB1004.ILE1616.net01342 ));
  inv_8_UCCLAB \ILAB1004.ILE1616.I666  ( .a(\ILAB1004.ILE1616.net01342 ), .x(\LLL15_PLL1<0> ));
  buftd4_UCCLAB \ILAB1004.I178  ( .a(\LLL15_PLL1<0> ), .en(VDD), .x(\ILAB1004.net015238 ));
  mux2p_2_UCCLAB \ILAB1004.I5605.I2  ( .d0(GND), .d1(\ILAB1004.net015238 ), .s0(VDD), .x(\ILAB1004.I5605.net33 ));
  invd16_seth_UCCLAB \ILAB1004.I5605.I3  ( .a(\ILAB1004.I5605.net33 ), .c(VDD), .x(\ILAB1004.Clk_int<2> ));
  mux2p_2_UCCLAB \ILAB1004.I5366.I82  ( .d0(GND), .d1(\ILAB1004.Clk_int<2> ), .s0(VDD), .x(\ILAB1004.I5366.net0119 ));
  invtd56_clk_UCCLAB \ILAB1004.I5366.I6  ( .a(\ILAB1004.I5366.net0119 ), .en(VDD), .x(\net16523<1> ));
  invtd56_UCCLAB \I3706.I4  ( .a(\net16523<1> ), .en(VDD), .x(\net10305<1> ));
  mux2_1_clk_P_UCCLAB \I3590.I17  ( .d0(\net10305<1> ), .d1(GND), .sl0(GND), .x(\I3590.net066 ));
  mux4p_0_UCCLAB \I3590.I13  ( .d0(GND), .d1(GND), .d2(GND), .d3(\I3590.net066 ), .sl0(VDD), .sl1(VDD), .x(\I3590.net78 ));
  invtd56_pd_clk_UCCLAB \I3590.I5  ( .a(\I3590.net78 ), .en(VDD), .x(\net10262<1> ));
  mux2p_2_UCCLAB \I3688.I4  ( .d0(\net10262<1> ), .d1(GND), .s0(GND), .x(\I3688.net43 ));
  invtd56_pd_clk_UCCLAB \I3688.I5  ( .a(\I3688.net43 ), .en(VDD), .x(\net10244<1> ));
  invtd56_pd_clk_UCCLAB \I3642.I2  ( .a(\net10244<1> ), .en(VDD), .x(\GCLK_s4<2> ));
  nand2_1_UCCLAB \ILAB0605.I5366.I72  ( .a(VDD), .b(\GCLK_s4<2> ), .x(\ILAB0605.I5366.net68 ));
  mux2d1i_1_P_UCCLAB \ILAB0605.I5366.I80  ( .d0(GND), .d1i(\ILAB0605.I5366.net68 ), .sl0(VDD), .x(\ILAB0605.I5366.net0106 ));
  invd52_UCCLAB \ILAB0605.I5366.I76  ( .a(\ILAB0605.I5366.net0106 ), .x(\ILAB0605.net15299<1> ));
  invd32_UCCLAB \ILAB0605.I5591.I1  ( .a(\ILAB0605.net15299<1> ), .x(\ILAB0605.Clk_LAB<2> ));
  mux2i_P_UCCLAB \IIO21.I0.I25  ( .d0(\IIO21.I0.net209 ), .d1(GND), .sl0(GND), .x(\IIO21.I0.net0153 ));
  invtd52_AVDD \IIO21.I0.I26  ( .a(\IIO21.I0.net0153 ), .en(VDD), .x(\LongBus_50<15> ));
  buftd52_UCCLAB \ILAB0506.I4801.I28  ( .a(\LongBus_50<15> ), .en(VDD), .x(\net8281<0> ));
  inv_4_UCCLAB \ILAB0506.ILE1606.I712  ( .a(\LongBus_50<15> ), .x(\ILAB0506.ILE1606.net0562 ));
  inv_4_UCCLAB \ILAB0606.ILE1016.I715  ( .a(\net8281<0> ), .x(\ILAB0606.ILE1016.net01339 ));
  inv_8_UCCLAB \ILAB0506.ILE1606.I666  ( .a(\ILAB0506.ILE1606.net0562 ), .x(\ILAB0506.net15881 ));
  buftd52_UCCLAB \ILAB0507.I4801.I28  ( .a(\LongBus_50<15> ), .en(VDD), .x(\net8302<0> ));
  buftd52_UCCLAB \ILAB0607.I4773.I29  ( .a(\net8302<0> ), .en(VDD), .x(\LongBus_49<15> ));
  inv_4_UCCLAB \ILAB0506.ILE1605.I710  ( .a(\LongBus_50<15> ), .x(\ILAB0506.ILE1605.net0558 ));
  inv_4_UCCLAB \ILAB0606.ILE0107.I713  ( .a(\LongBus_49<15> ), .x(\ILAB0606.ILE0107.net01342 ));
  inv_4_UCCLAB \ILAB0506.ILE0716.I714  ( .a(\net8281<0> ), .x(\ILAB0506.ILE0716.net01345 ));
  buftd4_UCCLAB \ILAB0506.I216  ( .a(\ILAB0506.net15881 ), .en(VDD), .x(\ILAB0506.net27188 ));
  mux2p_2_UCCLAB \ILAB0506.I5605.I0  ( .d0(\ILAB0506.net27188 ), .d1(GND), .s0(GND), .x(\ILAB0506.I5605.net29 ));
  invd16_seth_UCCLAB \ILAB0506.I5605.I1  ( .a(\ILAB0506.I5605.net29 ), .c(VDD), .x(\ILAB0506.Clk_int<3> ));
  mux2d1i_1_P_UCCLAB \ILAB0506.I5366.I81  ( .d0(\ILAB0506.Clk_int<3> ), .d1i(GND), .sl0(GND), .x(\ILAB0506.I5366.net0102 ));
  invd52_UCCLAB \ILAB0506.I5366.I77  ( .a(\ILAB0506.I5366.net0102 ), .x(\ILAB0506.net15299<0> ));
  invd32_UCCLAB \ILAB0506.I5591.I0  ( .a(\ILAB0506.net15299<0> ), .x(\ILAB0506.Clk_LAB<3> ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1615.Ivo1  ( .en(GND), .in(\ILAB0606.ILE1615.net2656 ), .out(\net14912<6> ));
  inv_8_UCCLAB \ILAB0606.ILE1615.I666  ( .a(\ILAB0606.ILE1615.net0541 ), .x(\ILAB0606.net22766 ));
  buf4_12_UCCLAB \ILAB0606.I4351  ( .a(\ILAB0606.net22766 ), .x(\ILAB0606.net39819 ));
  buftd52C_UCCLAB \ILAB0606.I4423  ( .a(\ILAB0606.net39819 ), .en(VDD), .x(\LongBus_48<15> ));
  buftd52_UCCLAB \ILAB0605.I4801.I28  ( .a(\LongBus_48<15> ), .en(VDD), .x(\net8290<0> ));
  buftd52C_UCCLAB \I1819.I28  ( .a(\net8290<0> ), .en(VDD), .x(\LongBus_33<15> ));
  buftd52_UCCLAB \ILAB1005.I4773.I29  ( .a(\LongBus_33<15> ), .en(VDD), .x(\LongBus_41<15> ));
  mux2i_P_UCCLAB \IIO26.I0.I16  ( .d0(GND), .d1(\LongBus_41<15> ), .sl0(VDD), .x(\IIO26.I0.net197 ));
  inv_8_UCCLAB \ILAB0606.ILE1415.I666  ( .a(\ILAB0606.ILE1415.net0541 ), .x(\ILAB0606.net19841 ));
  inv_8_UCCLAB \ILAB0606.ILE1416.I666  ( .a(\ILAB0606.net19841 ), .x(\net15029<1> ));
  buf4_12_UCCLAB \ILAB0606.I4369  ( .a(\net15029<1> ), .x(\ILAB0606.net27361 ));
  buftid52C_UCCLAB \ILAB0606.I4458  ( .a(\ILAB0606.net27361 ), .ne(GND), .x(\net8281<1> ));
  buftd52C_UCCLAB \I1823.I27  ( .a(\net8281<1> ), .en(VDD), .x(\LongBus_35<14> ));
  buftd52_UCCLAB \ILAB1006.I4773.I26  ( .a(\LongBus_35<14> ), .en(VDD), .x(\LongBus_41<14> ));
  mux2i_P_UCCLAB \IIO26.I1.I16  ( .d0(GND), .d1(\LongBus_41<14> ), .sl0(VDD), .x(\IIO26.I1.net197 ));
  inv_8_UCCLAB \ILAB0606.ILE1515.I666  ( .a(\ILAB0606.ILE1515.net0541 ), .x(\ILAB0606.net22046 ));
  inv_8_UCCLAB \ILAB0606.ILE1516.I666  ( .a(\ILAB0606.net22046 ), .x(\net15028<1> ));
  buf4_12_UCCLAB \ILAB0606.I4359  ( .a(\net15028<1> ), .x(\ILAB0606.net27381 ));
  buftid52C_UCCLAB \ILAB0606.I4460  ( .a(\ILAB0606.net27381 ), .ne(GND), .x(\net8281<2> ));
  buftd52C_UCCLAB \I1823.I31  ( .a(\net8281<2> ), .en(VDD), .x(\LongBus_35<13> ));
  buftd52_UCCLAB \ILAB1006.I4773.I30  ( .a(\LongBus_35<13> ), .en(VDD), .x(\LongBus_41<13> ));
  mux2i_P_UCCLAB \IIO26.I2.I16  ( .d0(GND), .d1(\LongBus_41<13> ), .sl0(VDD), .x(\IIO26.I2.net197 ));
  inv_8_UCCLAB \ILAB0706.ILE0113.I666  ( .a(\ILAB0706.ILE0113.net0541 ), .x(\ILAB0706.net21911 ));
  buf4_12_UCCLAB \ILAB0706.I4366  ( .a(\ILAB0706.net21911 ), .x(\ILAB0706.net38625 ));
  buftd52C_UCCLAB \ILAB0706.I4443  ( .a(\ILAB0706.net38625 ), .en(VDD), .x(\LongBus_47<4> ));
  buftd52_UCCLAB \ILAB0707.I4773.I40  ( .a(\LongBus_47<4> ), .en(VDD), .x(\net8302<11> ));
  buftd52C_UCCLAB \I1822.I40  ( .a(\net8302<11> ), .en(VDD), .x(\LongBus_37<4> ));
  buftd52_UCCLAB \ILAB1007.I4801.I41  ( .a(\LongBus_37<4> ), .en(VDD), .x(\LongBus_40<4> ));
  mux2i_P_UCCLAB \IIO26.I3.I16  ( .d0(\LongBus_40<4> ), .d1(GND), .sl0(GND), .x(\IIO26.I3.net197 ));
  inv_8_UCCLAB \ILAB0706.ILE0114.I666  ( .a(\ILAB0706.ILE0114.net0541 ), .x(\ILAB0706.net22271 ));
  buf4_12_UCCLAB \ILAB0706.I4387  ( .a(\ILAB0706.net22271 ), .x(\ILAB0706.net38763 ));
  buftd52C_UCCLAB \ILAB0706.I4445  ( .a(\ILAB0706.net38763 ), .en(VDD), .x(\LongBus_47<11> ));
  buftd52_UCCLAB \ILAB0707.I4773.I23  ( .a(\LongBus_47<11> ), .en(VDD), .x(\net8302<4> ));
  buftd52C_UCCLAB \I1822.I23  ( .a(\net8302<4> ), .en(VDD), .x(\LongBus_37<11> ));
  buftd52_UCCLAB \ILAB1007.I4773.I22  ( .a(\LongBus_37<11> ), .en(VDD), .x(\LongBus_41<11> ));
  mux2i_P_UCCLAB \IIO26.I4.I16  ( .d0(GND), .d1(\LongBus_41<11> ), .sl0(VDD), .x(\IIO26.I4.net197 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1313.Iho1  ( .en(GND), .in(\ILAB0606.ILE1313.net2656 ), .out(\net15072<0> ));
  inv_8_UCCLAB \ILAB0606.ILE1316.I666  ( .a(\net15072<0> ), .x(\net15030<1> ));
  buf4_12_UCCLAB \ILAB0606.I4396  ( .a(\net15030<1> ), .x(\ILAB0606.net27307 ));
  buftid52C_UCCLAB \ILAB0606.I4463  ( .a(\ILAB0606.net27307 ), .ne(GND), .x(\net8281<5> ));
  buftd52C_UCCLAB \I1823.I24  ( .a(\net8281<5> ), .en(VDD), .x(\LongBus_35<10> ));
  buftd52_UCCLAB \ILAB1006.I4773.I25  ( .a(\LongBus_35<10> ), .en(VDD), .x(\LongBus_41<10> ));
  mux2i_P_UCCLAB \IIO26.I5.I16  ( .d0(GND), .d1(\LongBus_41<10> ), .sl0(VDD), .x(\IIO26.I5.net197 ));
  inv_8_UCCLAB \ILAB0606.ILE1611.I666  ( .a(\ILAB0606.ILE1611.net0541 ), .x(\ILAB0606.net24386 ));
  buf4_12_UCCLAB \ILAB0606.I4399  ( .a(\ILAB0606.net24386 ), .x(\ILAB0606.net38760 ));
  buftd52C_UCCLAB \ILAB0606.I4451  ( .a(\ILAB0606.net38760 ), .en(VDD), .x(\LongBus_48<9> ));
  buftd52_UCCLAB \ILAB0605.I4801.I20  ( .a(\LongBus_48<9> ), .en(VDD), .x(\net8290<6> ));
  buftd52C_UCCLAB \I1819.I20  ( .a(\net8290<6> ), .en(VDD), .x(\LongBus_33<9> ));
  buftd52_UCCLAB \ILAB1005.I4773.I21  ( .a(\LongBus_33<9> ), .en(VDD), .x(\LongBus_41<9> ));
  mux2i_P_UCCLAB \IIO26.I6.I16  ( .d0(GND), .d1(\LongBus_41<9> ), .sl0(VDD), .x(\IIO26.I6.net197 ));
  inv_8_UCCLAB \ILAB0706.ILE0115.I666  ( .a(\ILAB0706.ILE0115.net0541 ), .x(\ILAB0706.net23666 ));
  buf4_12_UCCLAB \ILAB0706.I4370  ( .a(\ILAB0706.net23666 ), .x(\ILAB0706.net38388 ));
  buftd52C_UCCLAB \ILAB0706.I4435  ( .a(\ILAB0706.net38388 ), .en(VDD), .x(\LongBus_47<0> ));
  buftd52_UCCLAB \ILAB0707.I4773.I1  ( .a(\LongBus_47<0> ), .en(VDD), .x(\net8302<15> ));
  buftd52C_UCCLAB \I1822.I1  ( .a(\net8302<15> ), .en(VDD), .x(\LongBus_37<0> ));
  buftd52_UCCLAB \ILAB1007.I4801.I62895  ( .a(\LongBus_37<0> ), .en(VDD), .x(\LongBus_40<0> ));
  mux2i_P_UCCLAB \IIO26.I7.I16  ( .d0(\LongBus_40<0> ), .d1(GND), .sl0(GND), .x(\IIO26.I7.net197 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1114.Ihi7  ( .en(GND), .in(\ILAB0506.ILE1114.net2656 ), .out(\ILAB0506.net24952 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1114.Ivi5  ( .en(GND), .in(\ILAB0506.ILE1114.net2656 ), .out(\ILAB0506.net23537 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1114.Iho1  ( .en(GND), .in(\ILAB0506.ILE1114.net2656 ), .out(\net14778<1> ));
  inv_8_UCCLAB \ILAB0506.ILE1116.I666  ( .a(\net14778<1> ), .x(\net14730<1> ));
  buf4_12_UCCLAB \ILAB0506.I4408  ( .a(\net14730<1> ), .x(\ILAB0506.net27283 ));
  buftid52C_UCCLAB \ILAB0506.I4464  ( .a(\ILAB0506.net27283 ), .ne(GND), .x(\net8281<9> ));
  buftd52C_UCCLAB \I3749.I34  ( .a(\net8281<9> ), .en(VDD), .x(\LongBus_64<6> ));
  buftd52_UCCLAB \ILAB0306.I4801.I34  ( .a(\LongBus_64<6> ), .en(VDD), .x(\LongBus_54<6> ));
  mux2i_P_UCCLAB \IIO19.I1.I16  ( .d0(\LongBus_54<6> ), .d1(GND), .sl0(GND), .x(\IIO19.I1.net197 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE0912.Iho1  ( .en(GND), .in(\ILAB0506.ILE0912.net2656 ), .out(\ILAB0506.net18922 ));
  inv_8_UCCLAB \ILAB0506.ILE0912.I666  ( .a(\ILAB0506.ILE0912.net0541 ), .x(\ILAB0506.net18986 ));
  inv_4_UCCLAB \ILAB0506.ILE1013.I714  ( .a(\ILAB0506.net18986 ), .x(\ILAB0506.ILE1013.net01345 ));
  inv_8_UCCLAB \ILAB0506.ILE0916.I666  ( .a(\ILAB0506.net18922 ), .x(\net14732<1> ));
  buf4_12_UCCLAB \ILAB0506.I4401  ( .a(\net14732<1> ), .x(\ILAB0506.net27297 ));
  buftid52C_UCCLAB \ILAB0506.I4432  ( .a(\ILAB0506.net27297 ), .ne(GND), .x(\net8281<11> ));
  buftd52C_UCCLAB \I3749.I41  ( .a(\net8281<11> ), .en(VDD), .x(\LongBus_64<4> ));
  buftd52_UCCLAB \ILAB0306.I4801.I41  ( .a(\LongBus_64<4> ), .en(VDD), .x(\LongBus_54<4> ));
  mux2i_P_UCCLAB \IIO19.I3.I16  ( .d0(\LongBus_54<4> ), .d1(GND), .sl0(GND), .x(\IIO19.I3.net197 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE0912.Ivo3  ( .en(GND), .in(\ILAB0506.ILE0912.net2656 ), .out(\ILAB0506.net21690 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE0714.Ivo1  ( .en(GND), .in(\ILAB0506.ILE0714.net2656 ), .out(\ILAB0506.net23539 ));
  inv_8_UCCLAB \ILAB0506.ILE0714.I666  ( .a(\ILAB0506.ILE0714.net0541 ), .x(\ILAB0506.net19976 ));
  inv_4_UCCLAB \ILAB0506.ILE0813.I714  ( .a(\ILAB0506.net19976 ), .x(\ILAB0506.ILE0813.net01345 ));
  inv_4_UCCLAB \ILAB0506.ILE0613.I712  ( .a(\ILAB0506.net19976 ), .x(\ILAB0506.ILE0613.net0562 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE0714.Iho1  ( .en(GND), .in(\ILAB0506.ILE0714.net2656 ), .out(\net14794<1> ));
  inv_8_UCCLAB \ILAB0507.ILE0701.I666  ( .a(\net14794<1> ), .x(\net14734<0> ));
  buf4_12_UCCLAB \ILAB0507.I4395  ( .a(\net14734<0> ), .x(\ILAB0507.net39618 ));
  buftid52C_UCCLAB \ILAB0507.I4472  ( .a(\ILAB0507.net39618 ), .ne(GND), .x(\net8308<5> ));
  buftd52C_UCCLAB \I3752.I25  ( .a(\net8308<5> ), .en(VDD), .x(\LongBus_63<10> ));
  buftd52_UCCLAB \ILAB0307.I4772.I25  ( .a(\LongBus_63<10> ), .en(VDD), .x(\LongBus_55<10> ));
  mux2i_P_UCCLAB \IIO19.I5.I16  ( .d0(GND), .d1(\LongBus_55<10> ), .sl0(VDD), .x(\IIO19.I5.net197 ));
  inv_8_UCCLAB \ILAB0506.ILE0611.I666  ( .a(\ILAB0506.ILE0611.net0541 ), .x(\ILAB0506.net24116 ));
  inv_4_UCCLAB \ILAB0506.ILE0712.I714  ( .a(\ILAB0506.net24116 ), .x(\ILAB0506.ILE0712.net01345 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE0611.Ihi6  ( .en(GND), .in(\ILAB0506.ILE0611.net2656 ), .out(\ILAB0506.net19597 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE0612.Iho1  ( .en(GND), .in(\ILAB0506.net19597 ), .out(\ILAB0506.net19687 ));
  inv_8_UCCLAB \ILAB0506.ILE0616.I666  ( .a(\ILAB0506.net19687 ), .x(\net14735<1> ));
  buf4_12_UCCLAB \ILAB0506.I4405  ( .a(\net14735<1> ), .x(\ILAB0506.net27289 ));
  buftid52C_UCCLAB \ILAB0506.I4421  ( .a(\ILAB0506.net27289 ), .ne(GND), .x(\net8281<15> ));
  buftd52C_UCCLAB \I3749.I62895  ( .a(\net8281<15> ), .en(VDD), .x(\LongBus_64<0> ));
  buftd52_UCCLAB \ILAB0306.I4801.I62895  ( .a(\LongBus_64<0> ), .en(VDD), .x(\LongBus_54<0> ));
  mux2i_P_UCCLAB \IIO19.I7.I16  ( .d0(\LongBus_54<0> ), .d1(GND), .sl0(GND), .x(\IIO19.I7.net197 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE0511.Ivi7  ( .en(GND), .in(\ILAB0506.ILE0511.net2656 ), .out(\ILAB0506.net20389 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE0511.Ivi6  ( .en(GND), .in(\ILAB0506.ILE0511.net2656 ), .out(\ILAB0506.net21469 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE0511.Ivi5  ( .en(GND), .in(\ILAB0506.ILE0511.net2656 ), .out(\ILAB0506.net20387 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE0211.Ivi7  ( .en(GND), .in(\ILAB0506.net21469 ), .out(\net14777<1> ));
  inv_8_UCCLAB \ILAB0406.ILE1611.I666  ( .a(\net14777<1> ), .x(\ILAB0406.net24386 ));
  buf4_12_UCCLAB \ILAB0406.I4399  ( .a(\ILAB0406.net24386 ), .x(\ILAB0406.net38760 ));
  buftd52C_UCCLAB \ILAB0406.I4452  ( .a(\ILAB0406.net38760 ), .en(VDD), .x(\LongBus_52<14> ));
  buftd52_UCCLAB \ILAB0407.I4775.I27  ( .a(\LongBus_52<14> ), .en(VDD), .x(\net8308<1> ));
  buftd52C_UCCLAB \I3752.I26  ( .a(\net8308<1> ), .en(VDD), .x(\LongBus_63<14> ));
  buftd52_UCCLAB \ILAB0207.I4772.I26  ( .a(\LongBus_63<14> ), .en(VDD), .x(\LongBus_57<14> ));
  mux2i_P_UCCLAB \IIO18.I1.I16  ( .d0(GND), .d1(\LongBus_57<14> ), .sl0(VDD), .x(\IIO18.I1.net197 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE0512.Ivi7  ( .en(GND), .in(\ILAB0506.ILE0512.net2656 ), .out(\ILAB0506.net19084 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE0512.Ivi5  ( .en(GND), .in(\ILAB0506.ILE0512.net2656 ), .out(\ILAB0506.net19082 ));
  inv_8_UCCLAB \ILAB0506.ILE0316.I666  ( .a(\ILAB0506.net19082 ), .x(\net14738<1> ));
  buf4_12_UCCLAB \ILAB0506.I4398  ( .a(\net14738<1> ), .x(\ILAB0506.net27303 ));
  buftid52C_UCCLAB \ILAB0506.I4459  ( .a(\ILAB0506.net27303 ), .ne(GND), .x(\net8281<3> ));
  buftd52C_UCCLAB \I3749.I33  ( .a(\net8281<3> ), .en(VDD), .x(\LongBus_64<12> ));
  buftd52_UCCLAB \ILAB0206.I4773.I33  ( .a(\LongBus_64<12> ), .en(VDD), .x(\LongBus_57<12> ));
  mux2i_P_UCCLAB \IIO18.I3.I16  ( .d0(GND), .d1(\LongBus_57<12> ), .sl0(VDD), .x(\IIO18.I3.net197 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE0514.Ivi7  ( .en(GND), .in(\ILAB0506.ILE0514.net2656 ), .out(\ILAB0506.net19804 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE0514.Iho1  ( .en(GND), .in(\ILAB0506.ILE0514.net2656 ), .out(\net14802<1> ));
  inv_8_UCCLAB \ILAB0506.ILE0514.I666  ( .a(\ILAB0506.ILE0514.net0541 ), .x(\ILAB0506.net18311 ));
  inv_4_UCCLAB \ILAB0506.ILE0415.I712  ( .a(\ILAB0506.net18311 ), .x(\ILAB0506.ILE0415.net0562 ));
  inv_8_UCCLAB \ILAB0506.ILE0516.I666  ( .a(\net14802<1> ), .x(\net14736<1> ));
  buf4_12_UCCLAB \ILAB0506.I4380  ( .a(\net14736<1> ), .x(\ILAB0506.net27339 ));
  buftid52C_UCCLAB \ILAB0506.I4431  ( .a(\ILAB0506.net27339 ), .ne(GND), .x(\net8281<13> ));
  buftd52C_UCCLAB \I3749.I7  ( .a(\net8281<13> ), .en(VDD), .x(\LongBus_64<2> ));
  buftd52_UCCLAB \ILAB0206.I4801.I7  ( .a(\LongBus_64<2> ), .en(VDD), .x(\LongBus_56<2> ));
  mux2i_P_UCCLAB \IIO18.I5.I16  ( .d0(\LongBus_56<2> ), .d1(GND), .sl0(GND), .x(\IIO18.I5.net197 ));
  inv_8_UCCLAB \ILAB0506.ILE0614.I666  ( .a(\ILAB0506.ILE0614.net0541 ), .x(\ILAB0506.net19346 ));
  inv_4_UCCLAB \ILAB0506.ILE0515.I712  ( .a(\ILAB0506.net19346 ), .x(\ILAB0506.ILE0515.net0562 ));
  inv_4_UCCLAB \ILAB0506.ILE0515.I710  ( .a(\ILAB0506.net19346 ), .x(\ILAB0506.ILE0515.net0558 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE0614.Ivi7  ( .en(GND), .in(\ILAB0506.ILE0614.net2656 ), .out(\ILAB0506.net22144 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE0214.Ivi7  ( .en(GND), .in(\ILAB0506.net22144 ), .out(\net14765<1> ));
  inv_8_UCCLAB \ILAB0406.ILE1614.I666  ( .a(\net14765<1> ), .x(\ILAB0406.net20066 ));
  buf4_12_UCCLAB \ILAB0406.I4389  ( .a(\ILAB0406.net20066 ), .x(\ILAB0406.net37986 ));
  buftd52C_UCCLAB \ILAB0406.I4430  ( .a(\ILAB0406.net37986 ), .en(VDD), .x(\LongBus_52<0> ));
  buftd52_UCCLAB \ILAB0406.I4775.I1  ( .a(\LongBus_52<0> ), .en(VDD), .x(\net8314<15> ));
  buftd52C_UCCLAB \I3750.I62895  ( .a(\net8314<15> ), .en(VDD), .x(\LongBus_65<0> ));
  buftd52_UCCLAB \ILAB0206.I4775.I62895  ( .a(\LongBus_65<0> ), .en(VDD), .x(\LongBus_56<0> ));
  mux2i_P_UCCLAB \IIO18.I7.I16  ( .d0(\LongBus_56<0> ), .d1(GND), .sl0(GND), .x(\IIO18.I7.net197 ));
  inv_8_UCCLAB \ILAB0506.ILE1604.I666  ( .a(\ILAB0506.ILE1604.net0541 ), .x(\ILAB0506.net15476 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1604.Ivi7  ( .en(GND), .in(\ILAB0506.ILE1604.net2656 ), .out(\ILAB0506.net25384 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1604.Ihi7  ( .en(GND), .in(\ILAB0506.ILE1604.net2656 ), .out(\net13701<6> ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1603.Iho2  ( .en(GND), .in(\net13701<6> ), .out(\ILAB0506.net15458 ));
  inv_4_UCCLAB \ILAB0606.ILE0103.I715  ( .a(\ILAB0506.net15476 ), .x(\ILAB0606.ILE0103.net01339 ));
  inv_4_UCCLAB \ILAB0506.ILE1503.I711  ( .a(\ILAB0506.net15476 ), .x(\ILAB0506.ILE1503.net0560 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1404.Ihi5  ( .en(GND), .in(\ILAB0506.ILE1404.net2656 ), .out(\ILAB0506.net26303 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1404.Ihi7  ( .en(GND), .in(\ILAB0506.ILE1404.net2656 ), .out(\net13709<6> ));
  inv_8_UCCLAB \ILAB0506.ILE1404.I666  ( .a(\ILAB0506.ILE1404.net0541 ), .x(\ILAB0506.net20021 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1403.Iho2  ( .en(GND), .in(\net13709<6> ), .out(\ILAB0506.net20003 ));
  inv_4_UCCLAB \ILAB0506.ILE1503.I714  ( .a(\ILAB0506.net20021 ), .x(\ILAB0506.ILE1503.net01345 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1404.Ivo2  ( .en(GND), .in(\ILAB0506.ILE1404.net2656 ), .out(\ILAB0506.net25382 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1603.Ivo3  ( .en(GND), .in(\ILAB0506.net20003 ), .out(\net15111<4> ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0103.Ihi7  ( .en(GND), .in(\ILAB0606.ILE0103.net2656 ), .out(\net14063<3> ));
  inv_8_UCCLAB \ILAB0605.ILE0215.I666  ( .a(\ILAB0605.ILE0215.net0541 ), .x(\ILAB0605.net23756 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0215.Ivi7  ( .en(GND), .in(\ILAB0605.ILE0215.net2656 ), .out(\net14006<1> ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0115.Ivo2  ( .en(GND), .in(\net14006<1> ), .out(\ILAB0605.net24842 ));
  inv_4_UCCLAB \ILAB0605.ILE0116.I712  ( .a(\ILAB0605.net23756 ), .x(\ILAB0605.ILE0116.net0562 ));
  inv_4_UCCLAB \ILAB0605.ILE0116.I710  ( .a(\ILAB0605.net23756 ), .x(\ILAB0605.ILE0116.net0558 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0215.Ivo2  ( .en(GND), .in(\ILAB0605.ILE0215.net2656 ), .out(\ILAB0605.net22367 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0415.Ivo3  ( .en(GND), .in(\ILAB0605.net22367 ), .out(\ILAB0605.net22455 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1502.Ihi7  ( .en(GND), .in(\ILAB0506.ILE1502.net2656 ), .out(\net13705<1> ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1502.Ihi5  ( .en(GND), .in(\ILAB0506.ILE1502.net2656 ), .out(\net13705<5> ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1501.Iho2  ( .en(GND), .in(\net13705<1> ), .out(\ILAB0506.net20858 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1502.Ivi6  ( .en(GND), .in(\ILAB0506.ILE1502.net2656 ), .out(\ILAB0506.net26509 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0101.Ihi7  ( .en(GND), .in(\ILAB0606.ILE0101.net2656 ), .out(\net14063<0> ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1312.Ivo1  ( .en(GND), .in(\ILAB0505.ILE1312.net2656 ), .out(\net14018<0> ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1312.Ivo2  ( .en(GND), .in(\ILAB0505.ILE1312.net2656 ), .out(\ILAB0505.net19667 ));
  inv_8_UCCLAB \ILAB0505.ILE1312.I666  ( .a(\ILAB0505.ILE1312.net0541 ), .x(\ILAB0505.net22226 ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1512.Ivo3  ( .en(GND), .in(\ILAB0505.net19667 ), .out(\ILAB0505.net20115 ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1612.Ivo2  ( .en(GND), .in(\net14018<0> ), .out(\net14018<5> ));
  inv_4_UCCLAB \ILAB0505.ILE1411.I714  ( .a(\ILAB0505.net22226 ), .x(\ILAB0505.ILE1411.net01345 ));
  inv_4_UCCLAB \ILAB0505.ILE1413.I714  ( .a(\ILAB0505.net22226 ), .x(\ILAB0505.ILE1413.net01345 ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1610.Iho1  ( .en(GND), .in(\ILAB0505.ILE1610.net2656 ), .out(\ILAB0505.net24367 ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1610.Ivo1  ( .en(GND), .in(\ILAB0505.ILE1610.net2656 ), .out(\net14026<6> ));
  inv_8_UCCLAB \ILAB0505.ILE1610.I666  ( .a(\ILAB0505.ILE1610.net0541 ), .x(\ILAB0505.net16016 ));
  buftd4_UCCLAB \ILAB0505.I202  ( .a(\ILAB0505.net16016 ), .en(VDD), .x(\ILAB0505.net015238 ));
  mux2p_2_UCCLAB \ILAB0505.I5605.I2  ( .d0(GND), .d1(\ILAB0505.net015238 ), .s0(VDD), .x(\ILAB0505.I5605.net33 ));
  invd16_seth_UCCLAB \ILAB0505.I5605.I3  ( .a(\ILAB0505.I5605.net33 ), .c(VDD), .x(\ILAB0505.Clk_int<2> ));
  mux2d1i_1_P_UCCLAB \ILAB0505.I5366.I80  ( .d0(\ILAB0505.Clk_int<2> ), .d1i(GND), .sl0(GND), .x(\ILAB0505.I5366.net0106 ));
  invd52_UCCLAB \ILAB0505.I5366.I76  ( .a(\ILAB0505.I5366.net0106 ), .x(\ILAB0505.net15299<1> ));
  invd32_UCCLAB \ILAB0505.I5591.I1  ( .a(\ILAB0505.net15299<1> ), .x(\ILAB0505.Clk_LAB<2> ));
  inv_4_UCCLAB \ILAB0605.ILE0111.I714  ( .a(\ILAB0505.net16016 ), .x(\ILAB0605.ILE0111.net01345 ));
  inv_8_UCCLAB \ILAB0505.ILE1613.I666  ( .a(\ILAB0505.ILE1613.net0541 ), .x(\ILAB0505.net20111 ));
  buftd4_UCCLAB \ILAB0505.I189  ( .a(\ILAB0505.net20111 ), .en(VDD), .x(\ILAB0505.net27185 ));
  mux2p_2_UCCLAB \ILAB0505.I5605.I7  ( .d0(GND), .d1(\ILAB0505.net27185 ), .s0(VDD), .x(\ILAB0505.I5605.net21 ));
  invd16_seth_UCCLAB \ILAB0505.I5605.I6  ( .a(\ILAB0505.I5605.net21 ), .c(VDD), .x(\ILAB0505.Clk_int<0> ));
  mux2d1i_1_P_UCCLAB \ILAB0505.I5366.I78  ( .d0(\ILAB0505.Clk_int<0> ), .d1i(GND), .sl0(GND), .x(\ILAB0505.I5366.net0114 ));
  invd52_UCCLAB \ILAB0505.I5366.I74  ( .a(\ILAB0505.I5366.net0114 ), .x(\ILAB0505.net15299<3> ));
  invd32_UCCLAB \ILAB0505.I5591.I3  ( .a(\ILAB0505.net15299<3> ), .x(\ILAB0505.Clk_LAB<0> ));
  buf4_12_UCCLAB \ILAB0505.I4385  ( .a(\ILAB0505.net20111 ), .x(\ILAB0505.net38886 ));
  buftd52C_UCCLAB \ILAB0505.I4415  ( .a(\ILAB0505.net38886 ), .en(VDD), .x(\LongBus_50<4> ));
  buftd52_UCCLAB \ILAB0506.I4775.I40  ( .a(\LongBus_50<4> ), .en(VDD), .x(\net8314<11> ));
  inv_4_UCCLAB \ILAB0606.ILE0301.I713  ( .a(\net8314<11> ), .x(\ILAB0606.ILE0301.net01342 ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1214.Ivo2  ( .en(GND), .in(\ILAB0505.ILE1214.net2656 ), .out(\ILAB0505.net19847 ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1214.Iho2  ( .en(GND), .in(\ILAB0505.ILE1214.net2656 ), .out(\ILAB0505.net23423 ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1414.Ivo3  ( .en(GND), .in(\ILAB0505.net19847 ), .out(\ILAB0505.net22050 ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1216.Iho3  ( .en(GND), .in(\ILAB0505.net23423 ), .out(\net13717<4> ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1214.Ivi6  ( .en(GND), .in(\ILAB0505.ILE1214.net2656 ), .out(\ILAB0505.net23269 ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1314.Ivo1  ( .en(GND), .in(\ILAB0505.net23269 ), .out(\net14010<0> ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0114.Ivo1  ( .en(GND), .in(\net14010<0> ), .out(\ILAB0605.net19804 ));
  inv_8_UCCLAB \ILAB0505.ILE1314.I666  ( .a(\ILAB0505.ILE1314.net0541 ), .x(\ILAB0505.net21011 ));
  inv_4_UCCLAB \ILAB0505.ILE1413.I715  ( .a(\ILAB0505.net21011 ), .x(\ILAB0505.ILE1413.net01339 ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1314.Ivo2  ( .en(GND), .in(\ILAB0505.ILE1314.net2656 ), .out(\ILAB0505.net22052 ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1414.Ivo1  ( .en(GND), .in(\ILAB0505.ILE1414.net2656 ), .out(\net14010<1> ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0613.Ihi6  ( .en(GND), .in(\ILAB0605.ILE0613.net2656 ), .out(\ILAB0605.net24097 ));
  inv_8_UCCLAB \ILAB0605.ILE0613.I666  ( .a(\ILAB0605.ILE0613.net0541 ), .x(\ILAB0605.net19706 ));
  inv_4_UCCLAB \ILAB0605.ILE0514.I710  ( .a(\ILAB0605.net19706 ), .x(\ILAB0605.ILE0514.net0558 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0613.Ivi5  ( .en(GND), .in(\ILAB0605.ILE0613.net2656 ), .out(\ILAB0605.net19352 ));
  inv_8_UCCLAB \ILAB0605.ILE0515.I666  ( .a(\ILAB0605.ILE0515.net0541 ), .x(\ILAB0605.net19796 ));
  inv_4_UCCLAB \ILAB0605.ILE0416.I712  ( .a(\ILAB0605.net19796 ), .x(\ILAB0605.ILE0416.net0562 ));
  inv_4_UCCLAB \ILAB0605.ILE0414.I712  ( .a(\ILAB0605.net19796 ), .x(\ILAB0605.ILE0414.net0562 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0515.Iho1  ( .en(GND), .in(\ILAB0605.ILE0515.net2656 ), .out(\net14047<3> ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0414.Ivi7  ( .en(GND), .in(\ILAB0605.ILE0414.net2656 ), .out(\net14010<6> ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0113.Ivo2  ( .en(GND), .in(\ILAB0605.ILE0113.net2656 ), .out(\ILAB0605.net23177 ));
  inv_8_UCCLAB \ILAB0605.ILE0113.I666  ( .a(\ILAB0605.ILE0113.net0541 ), .x(\ILAB0605.net21911 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0313.Ivo3  ( .en(GND), .in(\ILAB0605.net23177 ), .out(\ILAB0605.net26100 ));
  inv_4_UCCLAB \ILAB0605.ILE0212.I713  ( .a(\ILAB0605.net21911 ), .x(\ILAB0605.ILE0212.net01342 ));
  inv_4_UCCLAB \ILAB0605.ILE0214.I714  ( .a(\ILAB0605.net21911 ), .x(\ILAB0605.ILE0214.net01345 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0113.Ivo3  ( .en(GND), .in(\ILAB0605.ILE0113.net2656 ), .out(\ILAB0605.net23085 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0313.Iho1  ( .en(GND), .in(\ILAB0605.ILE0313.net2656 ), .out(\net14055<0> ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0313.Ivo1  ( .en(GND), .in(\ILAB0605.ILE0313.net2656 ), .out(\ILAB0605.net19984 ));
  inv_8_UCCLAB \ILAB0605.ILE0313.I666  ( .a(\ILAB0605.ILE0313.net0541 ), .x(\ILAB0605.net24926 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0316.Iho2  ( .en(GND), .in(\net14055<0> ), .out(\net14055<5> ));
  inv_4_UCCLAB \ILAB0605.ILE0412.I715  ( .a(\ILAB0605.net24926 ), .x(\ILAB0605.ILE0412.net01339 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0314.Ivi5  ( .en(GND), .in(\ILAB0605.ILE0314.net2656 ), .out(\ILAB0605.net23807 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0114.Ihi6  ( .en(GND), .in(\ILAB0605.net23807 ), .out(\ILAB0605.net23197 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0114.Iho1  ( .en(GND), .in(\ILAB0605.ILE0114.net2656 ), .out(\net14063<1> ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0711.Ivi6  ( .en(GND), .in(\ILAB0605.ILE0711.net2656 ), .out(\ILAB0605.net18499 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0510.Iho3  ( .en(GND), .in(\ILAB0605.ILE0510.net2656 ), .out(\ILAB0605.net23919 ));
  inv_8_UCCLAB \ILAB0605.ILE0510.I666  ( .a(\ILAB0605.ILE0510.net0541 ), .x(\ILAB0605.net19121 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0510.Ivi5  ( .en(GND), .in(\ILAB0605.ILE0510.net2656 ), .out(\ILAB0605.net23942 ));
  inv_4_UCCLAB \ILAB0605.ILE0411.I712  ( .a(\ILAB0605.net19121 ), .x(\ILAB0605.ILE0411.net0562 ));
  inv_4_UCCLAB \ILAB0605.ILE0611.I714  ( .a(\ILAB0605.net19121 ), .x(\ILAB0605.ILE0611.net01345 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0511.Iho3  ( .en(GND), .in(\ILAB0605.ILE0511.net2656 ), .out(\ILAB0605.net20364 ));
  inv_8_UCCLAB \ILAB0605.ILE0511.I666  ( .a(\ILAB0605.ILE0511.net0541 ), .x(\ILAB0605.net23936 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0511.Ivi7  ( .en(GND), .in(\ILAB0605.ILE0511.net2656 ), .out(\ILAB0605.net20389 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0411.Ivo2  ( .en(GND), .in(\ILAB0605.net20389 ), .out(\ILAB0605.net21467 ));
  inv_4_UCCLAB \ILAB0605.ILE0412.I712  ( .a(\ILAB0605.net23936 ), .x(\ILAB0605.ILE0412.net0562 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0215.Iho2  ( .en(GND), .in(\ILAB0605.net20364 ), .out(\net14059<2> ));
  inv_8_UCCLAB \ILAB0506.ILE1202.I666  ( .a(\ILAB0506.ILE1202.net0541 ), .x(\ILAB0506.net15521 ));
  inv_4_UCCLAB \ILAB0506.ILE1301.I715  ( .a(\ILAB0506.net15521 ), .x(\ILAB0506.ILE1301.net01339 ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1115.Ivo2  ( .en(GND), .in(\ILAB0505.ILE1115.net2656 ), .out(\ILAB0505.net24302 ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1315.Ivo3  ( .en(GND), .in(\ILAB0505.net24302 ), .out(\ILAB0505.net22725 ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1115.Ivo3  ( .en(GND), .in(\ILAB0505.ILE1115.net2656 ), .out(\ILAB0505.net24435 ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1115.Iho2  ( .en(GND), .in(\ILAB0505.ILE1115.net2656 ), .out(\net13721<2> ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1101.Iho3  ( .en(GND), .in(\net13721<2> ), .out(\ILAB0506.net16584 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1301.Ivo1  ( .en(GND), .in(\ILAB0506.ILE1301.net2656 ), .out(\net15119<0> ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1601.Ivo2  ( .en(GND), .in(\net15119<0> ), .out(\net15119<5> ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1301.Ivi6  ( .en(GND), .in(\ILAB0506.ILE1301.net2656 ), .out(\ILAB0506.net20839 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1401.Ivo1  ( .en(GND), .in(\ILAB0506.net20839 ), .out(\net15119<1> ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0101.Ivo2  ( .en(GND), .in(\net15119<1> ), .out(\ILAB0606.net17867 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0301.Ivo3  ( .en(GND), .in(\ILAB0606.net17867 ), .out(\ILAB0606.net20745 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0106.Ihi5  ( .en(GND), .in(\ILAB0606.ILE0106.net2656 ), .out(\ILAB0606.net22928 ));
  inv_8_UCCLAB \ILAB0606.ILE0106.I666  ( .a(\ILAB0606.ILE0106.net0541 ), .x(\ILAB0606.net19751 ));
  inv_4_UCCLAB \ILAB0606.ILE0205.I713  ( .a(\ILAB0606.net19751 ), .x(\ILAB0606.ILE0205.net01342 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0104.Ivi6  ( .en(GND), .in(\ILAB0606.net22928 ), .out(\net15107<1> ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0207.Ihi7  ( .en(GND), .in(\ILAB0606.ILE0207.net2656 ), .out(\ILAB0606.net23827 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0207.Ivi7  ( .en(GND), .in(\ILAB0606.ILE0207.net2656 ), .out(\net15095<1> ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0207.Ihi6  ( .en(GND), .in(\ILAB0606.ILE0207.net2656 ), .out(\ILAB0606.net20227 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0204.Ivi5  ( .en(GND), .in(\ILAB0606.net20227 ), .out(\net15107<5> ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0104.Ihi7  ( .en(GND), .in(\ILAB0606.ILE0104.net2656 ), .out(\net14063<6> ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0104.Ihi6  ( .en(GND), .in(\ILAB0606.ILE0104.net2656 ), .out(\ILAB0606.net16717 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0201.Iho3  ( .en(GND), .in(\ILAB0606.ILE0201.net2656 ), .out(\ILAB0606.net16944 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0406.Ihi5  ( .en(GND), .in(\ILAB0606.ILE0406.net2656 ), .out(\ILAB0606.net15548 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0406.Ivi7  ( .en(GND), .in(\ILAB0606.ILE0406.net2656 ), .out(\net15099<6> ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0406.Ihi6  ( .en(GND), .in(\ILAB0606.ILE0406.net2656 ), .out(\ILAB0606.net20182 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0403.Ihi7  ( .en(GND), .in(\ILAB0606.net20182 ), .out(\net14051<3> ));
  inv_8_UCCLAB \ILAB0606.ILE0306.I666  ( .a(\ILAB0606.ILE0306.net0541 ), .x(\ILAB0606.net23351 ));
  inv_4_UCCLAB \ILAB0606.ILE0205.I710  ( .a(\ILAB0606.net23351 ), .x(\ILAB0606.ILE0205.net0558 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0306.Ivi7  ( .en(GND), .in(\ILAB0606.ILE0306.net2656 ), .out(\net15099<3> ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0306.Ihi7  ( .en(GND), .in(\ILAB0606.ILE0306.net2656 ), .out(\ILAB0606.net26797 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0302.Ihi7  ( .en(GND), .in(\ILAB0606.net26797 ), .out(\net14055<1> ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0206.Ihi7  ( .en(GND), .in(\ILAB0606.ILE0206.net2656 ), .out(\ILAB0606.net26752 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0504.Ihi5  ( .en(GND), .in(\ILAB0606.ILE0504.net2656 ), .out(\ILAB0606.net26258 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0504.Ihi7  ( .en(GND), .in(\ILAB0606.ILE0504.net2656 ), .out(\net14047<6> ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0516.Ivi7  ( .en(GND), .in(\net14047<6> ), .out(\ILAB0605.net17014 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0504.Ivi5  ( .en(GND), .in(\ILAB0606.ILE0504.net2656 ), .out(\ILAB0606.net25022 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0304.Ivi6  ( .en(GND), .in(\ILAB0606.net25022 ), .out(\net15107<6> ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0402.Iho1  ( .en(GND), .in(\ILAB0606.ILE0402.net2656 ), .out(\ILAB0606.net26212 ));
  inv_8_UCCLAB \ILAB0606.ILE0402.I666  ( .a(\ILAB0606.ILE0402.net0541 ), .x(\ILAB0606.net20741 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0402.Ivi5  ( .en(GND), .in(\ILAB0606.ILE0402.net2656 ), .out(\ILAB0606.net26237 ));
  inv_4_UCCLAB \ILAB0606.ILE0301.I712  ( .a(\ILAB0606.net20741 ), .x(\ILAB0606.ILE0301.net0562 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0402.Iho3  ( .en(GND), .in(\ILAB0606.ILE0402.net2656 ), .out(\ILAB0606.net26214 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0204.Ihi7  ( .en(GND), .in(\ILAB0606.ILE0204.net2656 ), .out(\net14059<6> ));
  inv_8_UCCLAB \ILAB0505.ILE1415.I666  ( .a(\ILAB0505.ILE1415.net0541 ), .x(\ILAB0505.net19841 ));
  inv_4_UCCLAB \ILAB0505.ILE1514.I713  ( .a(\ILAB0505.net19841 ), .x(\ILAB0505.ILE1514.net01342 ));
  inv_4_UCCLAB \ILAB0505.ILE1516.I714  ( .a(\ILAB0505.net19841 ), .x(\ILAB0505.ILE1516.net01345 ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1415.Ivo3  ( .en(GND), .in(\ILAB0505.ILE1415.net2656 ), .out(\ILAB0505.net22815 ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1415.Ivo2  ( .en(GND), .in(\ILAB0505.ILE1415.net2656 ), .out(\ILAB0505.net24257 ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1511.Iho1  ( .en(GND), .in(\ILAB0505.ILE1511.net2656 ), .out(\ILAB0505.net21262 ));
  inv_8_UCCLAB \ILAB0505.ILE1511.I666  ( .a(\ILAB0505.ILE1511.net0541 ), .x(\ILAB0505.net24071 ));
  inv_4_UCCLAB \ILAB0505.ILE1612.I715  ( .a(\ILAB0505.net24071 ), .x(\ILAB0505.ILE1612.net01339 ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1511.Ivo3  ( .en(GND), .in(\ILAB0505.ILE1511.net2656 ), .out(\ILAB0505.net22005 ));
  inv_8_UCCLAB \ILAB0505.ILE1614.I666  ( .a(\ILAB0505.ILE1614.net0541 ), .x(\ILAB0505.net20066 ));
  buftd4_UCCLAB \ILAB0505.I183  ( .a(\ILAB0505.net20066 ), .en(VDD), .x(\ILAB0505.net27191 ));
  mux2p_2_UCCLAB \ILAB0505.I5605.I4  ( .d0(GND), .d1(\ILAB0505.net27191 ), .s0(VDD), .x(\ILAB0505.I5605.net25 ));
  invd16_seth_UCCLAB \ILAB0505.I5605.I5  ( .a(\ILAB0505.I5605.net25 ), .c(VDD), .x(\ILAB0505.Clk_int<1> ));
  mux2p_2_UCCLAB \ILAB0505.I5366.I83  ( .d0(\ILAB0505.Clk_int<1> ), .d1(GND), .s0(GND), .x(\ILAB0505.I5366.net0122 ));
  invtd56_clk_UCCLAB \ILAB0505.I5366.I8  ( .a(\ILAB0505.I5366.net0122 ), .en(VDD), .x(\net10221<0> ));
  invtd56_UCCLAB \I3697.I3  ( .a(\net10221<0> ), .en(VDD), .x(\net10247<0> ));
  mux2p_2_UCCLAB \I3688.I6  ( .d0(GND), .d1(\net10247<0> ), .s0(VDD), .x(\I3688.net47 ));
  invtd56_pd_clk_UCCLAB \I3688.I0  ( .a(\I3688.net47 ), .en(VDD), .x(\net10244<0> ));
  invtd56_pd_clk_UCCLAB \I3642.I1  ( .a(\net10244<0> ), .en(VDD), .x(\GCLK_s4<3> ));
  nand2_1_UCCLAB \ILAB0605.I5366.I73  ( .a(VDD), .b(\GCLK_s4<3> ), .x(\ILAB0605.I5366.net66 ));
  mux2d1i_1_P_UCCLAB \ILAB0605.I5366.I81  ( .d0(GND), .d1i(\ILAB0605.I5366.net66 ), .sl0(VDD), .x(\ILAB0605.I5366.net0102 ));
  invd52_UCCLAB \ILAB0605.I5366.I77  ( .a(\ILAB0605.I5366.net0102 ), .x(\ILAB0605.net15299<0> ));
  invd32_UCCLAB \ILAB0605.I5591.I0  ( .a(\ILAB0605.net15299<0> ), .x(\ILAB0605.Clk_LAB<3> ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0310.Iho3  ( .en(GND), .in(\ILAB0605.ILE0310.net2656 ), .out(\ILAB0605.net25899 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0310.Iho1  ( .en(GND), .in(\ILAB0605.ILE0310.net2656 ), .out(\ILAB0605.net25897 ));
  inv_8_UCCLAB \ILAB0605.ILE0310.I666  ( .a(\ILAB0605.ILE0310.net0541 ), .x(\ILAB0605.net16511 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0310.Ivi7  ( .en(GND), .in(\ILAB0605.ILE0310.net2656 ), .out(\net14026<3> ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0210.Ivo2  ( .en(GND), .in(\net14026<3> ), .out(\ILAB0605.net23897 ));
  inv_4_UCCLAB \ILAB0605.ILE0211.I712  ( .a(\ILAB0605.net16511 ), .x(\ILAB0605.ILE0211.net0562 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0313.Iho2  ( .en(GND), .in(\ILAB0605.net25897 ), .out(\ILAB0605.net23153 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0315.Iho3  ( .en(GND), .in(\ILAB0605.net23153 ), .out(\ILAB0605.net24819 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0212.Iho3  ( .en(GND), .in(\ILAB0605.net23897 ), .out(\ILAB0605.net22299 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0601.Ihi5  ( .en(GND), .in(\ILAB0606.ILE0601.net2656 ), .out(\net14043<2> ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0601.Ihi7  ( .en(GND), .in(\ILAB0606.ILE0601.net2656 ), .out(\net14043<0> ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0601.Ihi6  ( .en(GND), .in(\ILAB0606.ILE0601.net2656 ), .out(\net14043<1> ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0601.Ivi6  ( .en(GND), .in(\ILAB0606.ILE0601.net2656 ), .out(\ILAB0606.net20524 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0301.Ivi7  ( .en(GND), .in(\ILAB0606.net20524 ), .out(\net15119<3> ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0415.Ivi6  ( .en(GND), .in(\net14043<1> ), .out(\ILAB0605.net22459 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0315.Iho1  ( .en(GND), .in(\ILAB0605.ILE0315.net2656 ), .out(\net14055<3> ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0302.Iho2  ( .en(GND), .in(\net14055<3> ), .out(\ILAB0606.net26798 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0302.Ivi5  ( .en(GND), .in(\ILAB0606.net26798 ), .out(\ILAB0606.net26822 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0202.Ivi7  ( .en(GND), .in(\ILAB0606.ILE0202.net2656 ), .out(\net15115<1> ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0102.Iho1  ( .en(GND), .in(\ILAB0606.ILE0102.net2656 ), .out(\ILAB0606.net26707 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0102.Ivi7  ( .en(GND), .in(\ILAB0606.ILE0102.net2656 ), .out(\net15115<0> ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0106.Iho1  ( .en(GND), .in(\ILAB0606.net26707 ), .out(\ILAB0606.net17257 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0109.Iho2  ( .en(GND), .in(\ILAB0606.net17257 ), .out(\ILAB0606.net16403 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0111.Iho3  ( .en(GND), .in(\ILAB0606.net16403 ), .out(\ILAB0606.net23199 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1306.Iho1  ( .en(GND), .in(\net15115<0> ), .out(\ILAB0506.net18697 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1310.Iho1  ( .en(GND), .in(\ILAB0506.net18697 ), .out(\ILAB0506.net24682 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0511.Ivo1  ( .en(GND), .in(\ILAB0606.net23199 ), .out(\ILAB0606.net18994 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0811.Ivo2  ( .en(GND), .in(\ILAB0606.net18994 ), .out(\ILAB0606.net22682 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1011.Ivo3  ( .en(GND), .in(\ILAB0606.net22682 ), .out(\ILAB0606.net23040 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1305.Iho2  ( .en(GND), .in(\net15115<0> ), .out(\ILAB0506.net15908 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0301.Iho2  ( .en(GND), .in(\ILAB0606.ILE0301.net2656 ), .out(\ILAB0606.net17843 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0302.Iho3  ( .en(GND), .in(\ILAB0606.ILE0302.net2656 ), .out(\ILAB0606.net26799 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0214.Iho1  ( .en(GND), .in(\ILAB0605.ILE0214.net2656 ), .out(\net14059<1> ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0201.Iho2  ( .en(GND), .in(\net14059<1> ), .out(\ILAB0606.net16943 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0203.Ivo1  ( .en(GND), .in(\ILAB0606.ILE0203.net2656 ), .out(\ILAB0606.net17689 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0416.Ivi7  ( .en(GND), .in(\ILAB0605.ILE0416.net2656 ), .out(\net14002<6> ));
  inv_8_UCCLAB \ILAB0506.ILE1602.I666  ( .a(\ILAB0506.ILE1602.net0541 ), .x(\ILAB0506.net20561 ));
  buftd4_UCCLAB \ILAB0506.I233  ( .a(\ILAB0506.net20561 ), .en(VDD), .x(\ILAB0506.net027160 ));
  mux2p_2_UCCLAB \ILAB0506.I5605.I7  ( .d0(\ILAB0506.net027160 ), .d1(GND), .s0(GND), .x(\ILAB0506.I5605.net21 ));
  invd16_seth_UCCLAB \ILAB0506.I5605.I6  ( .a(\ILAB0506.I5605.net21 ), .c(VDD), .x(\ILAB0506.Clk_int<0> ));
  mux2p_2_UCCLAB \ILAB0506.I5366.I82  ( .d0(\ILAB0506.Clk_int<0> ), .d1(GND), .s0(GND), .x(\ILAB0506.I5366.net0119 ));
  invtd56_clk_UCCLAB \ILAB0506.I5366.I6  ( .a(\ILAB0506.I5366.net0119 ), .en(VDD), .x(\net10221<1> ));
  invtd56_UCCLAB \I3697.I4  ( .a(\net10221<1> ), .en(VDD), .x(\net10247<1> ));
  mux2p_2_UCCLAB \I3688.I2  ( .d0(GND), .d1(\net10247<1> ), .s0(VDD), .x(\I3688.net35 ));
  invtd56_pd_clk_UCCLAB \I3688.I9  ( .a(\I3688.net35 ), .en(VDD), .x(\net10244<3> ));
  invtd56_pd_clk_UCCLAB \I3642.I4  ( .a(\net10244<3> ), .en(VDD), .x(\GCLK_s4<0> ));
  nand2_1_UCCLAB \ILAB0605.I5366.I0  ( .a(VDD), .b(\GCLK_s4<0> ), .x(\ILAB0605.I5366.net64 ));
  mux2d1i_1_P_UCCLAB \ILAB0605.I5366.I78  ( .d0(GND), .d1i(\ILAB0605.I5366.net64 ), .sl0(VDD), .x(\ILAB0605.I5366.net0114 ));
  invd52_UCCLAB \ILAB0605.I5366.I74  ( .a(\ILAB0605.I5366.net0114 ), .x(\ILAB0605.net15299<3> ));
  invd32_UCCLAB \ILAB0605.I5591.I3  ( .a(\ILAB0605.net15299<3> ), .x(\ILAB0605.Clk_LAB<0> ));
  inv_8_UCCLAB \ILAB0605.ILE0415.I666  ( .a(\ILAB0605.ILE0415.net0541 ), .x(\ILAB0605.net19256 ));
  inv_4_UCCLAB \ILAB0605.ILE0316.I711  ( .a(\ILAB0605.net19256 ), .x(\ILAB0605.ILE0316.net0560 ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1514.Ivo1  ( .en(GND), .in(\ILAB0505.ILE1514.net2656 ), .out(\net14010<3> ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0214.Ivo2  ( .en(GND), .in(\net14010<3> ), .out(\ILAB0605.net19262 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0216.Ivo1  ( .en(GND), .in(\ILAB0605.ILE0216.net2656 ), .out(\ILAB0605.net18859 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0316.Iho1  ( .en(GND), .in(\ILAB0605.ILE0316.net2656 ), .out(\net14055<6> ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0303.Ivi5  ( .en(GND), .in(\ILAB0606.ILE0303.net2656 ), .out(\ILAB0606.net23582 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0303.Iho1  ( .en(GND), .in(\ILAB0606.ILE0303.net2656 ), .out(\ILAB0606.net23557 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0306.Iho2  ( .en(GND), .in(\ILAB0606.net23557 ), .out(\ILAB0606.net17528 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0303.Ivi6  ( .en(GND), .in(\ILAB0606.ILE0303.net2656 ), .out(\net15111<6> ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0303.Ivo2  ( .en(GND), .in(\ILAB0606.ILE0303.net2656 ), .out(\ILAB0606.net20162 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0103.Ivi6  ( .en(GND), .in(\ILAB0606.net23582 ), .out(\net15111<1> ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0503.Ivo3  ( .en(GND), .in(\ILAB0606.net20162 ), .out(\ILAB0606.net17685 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0307.Iho1  ( .en(GND), .in(\ILAB0606.net23557 ), .out(\ILAB0606.net25852 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0310.Iho2  ( .en(GND), .in(\ILAB0606.net25852 ), .out(\ILAB0606.net25898 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0311.Iho1  ( .en(GND), .in(\ILAB0606.net25852 ), .out(\ILAB0606.net23377 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0312.Iho3  ( .en(GND), .in(\ILAB0606.net25898 ), .out(\ILAB0606.net24909 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0314.Iho2  ( .en(GND), .in(\ILAB0606.net23377 ), .out(\ILAB0606.net23783 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1403.Ivi7  ( .en(GND), .in(\net15111<1> ), .out(\ILAB0506.net20029 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0407.Ivo1  ( .en(GND), .in(\ILAB0606.net23557 ), .out(\ILAB0606.net25249 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0807.Ivo1  ( .en(GND), .in(\ILAB0606.net25249 ), .out(\ILAB0606.net17059 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1307.Ivi7  ( .en(GND), .in(\ILAB0606.net23582 ), .out(\ILAB0506.net17149 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1509.Ivi7  ( .en(GND), .in(\ILAB0606.net25852 ), .out(\ILAB0506.net18049 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0409.Ivo1  ( .en(GND), .in(\ILAB0606.net25852 ), .out(\ILAB0606.net17644 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1207.Ivo1  ( .en(GND), .in(\ILAB0606.net17059 ), .out(\ILAB0606.net15349 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0714.Ivo1  ( .en(GND), .in(\ILAB0606.net23783 ), .out(\ILAB0606.net23539 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0712.Ivo1  ( .en(GND), .in(\ILAB0606.net24909 ), .out(\ILAB0606.net21784 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0809.Ivo1  ( .en(GND), .in(\ILAB0606.net17644 ), .out(\ILAB0606.net16294 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1211.Iho1  ( .en(GND), .in(\ILAB0606.net15349 ), .out(\ILAB0606.net22567 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1007.Iho1  ( .en(GND), .in(\ILAB0506.net20029 ), .out(\ILAB0506.net25807 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE0911.Iho1  ( .en(GND), .in(\ILAB0506.net17149 ), .out(\ILAB0506.net18967 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1011.Iho1  ( .en(GND), .in(\ILAB0506.net25807 ), .out(\ILAB0506.net22657 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1405.Ihi7  ( .en(GND), .in(\ILAB0506.ILE1405.net2656 ), .out(\ILAB0506.net20812 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1405.Ivo1  ( .en(GND), .in(\ILAB0506.ILE1405.net2656 ), .out(\net15103<1> ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1401.Ihi7  ( .en(GND), .in(\ILAB0506.net20812 ), .out(\net13709<0> ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0105.Ivo2  ( .en(GND), .in(\net15103<1> ), .out(\ILAB0606.net23357 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1503.Ivo1  ( .en(GND), .in(\ILAB0506.net20812 ), .out(\net15111<3> ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1413.Ihi7  ( .en(GND), .in(\net13709<0> ), .out(\ILAB0505.net18067 ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1511.Ivo1  ( .en(GND), .in(\ILAB0505.net18067 ), .out(\net14022<3> ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0211.Ivo2  ( .en(GND), .in(\net14022<3> ), .out(\ILAB0605.net19892 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1405.Ivi5  ( .en(GND), .in(\ILAB0506.ILE1405.net2656 ), .out(\ILAB0506.net25067 ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1314.Ihi7  ( .en(GND), .in(\ILAB0506.net25067 ), .out(\ILAB0505.net24682 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0209.Ivo1  ( .en(GND), .in(\ILAB0505.net18067 ), .out(\ILAB0605.net15439 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0415.Ivo1  ( .en(GND), .in(\net15111<3> ), .out(\ILAB0605.net22099 ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1612.Ivo3  ( .en(GND), .in(\net13709<0> ), .out(\net14018<4> ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0609.Ivo1  ( .en(GND), .in(\ILAB0605.net15439 ), .out(\ILAB0605.net16339 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0213.Ivo1  ( .en(GND), .in(\net13709<0> ), .out(\ILAB0605.net19354 ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1512.Ivo1  ( .en(GND), .in(\ILAB0505.net18067 ), .out(\net14018<3> ));
  inv_8_UCCLAB \ILAB0505.ILE1416.I666  ( .a(\net13709<0> ), .x(\net13670<1> ));
  buf4_12_UCCLAB \ILAB0505.I4369  ( .a(\net13670<1> ), .x(\ILAB0505.net27361 ));
  buftid52C_UCCLAB \ILAB0505.I4466  ( .a(\ILAB0505.net27361 ), .ne(GND), .x(\net8290<14> ));
  inv_4_UCCLAB \ILAB0605.ILE0516.I713  ( .a(\net8290<14> ), .x(\ILAB0605.ILE0516.net01342 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0302.Ivo1  ( .en(GND), .in(\net15103<1> ), .out(\ILAB0606.net26464 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0107.Ivo1  ( .en(GND), .in(\ILAB0606.ILE0107.net2656 ), .out(\net15022<6> ));
  inv_8_UCCLAB \ILAB0606.ILE0105.I666  ( .a(\ILAB0606.ILE0105.net0541 ), .x(\ILAB0606.net22946 ));
  inv_4_UCCLAB \ILAB0506.ILE1606.I710  ( .a(\ILAB0606.net22946 ), .x(\ILAB0506.ILE1606.net0558 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1606.Ivo3  ( .en(GND), .in(\ILAB0506.ILE1606.net2656 ), .out(\net15099<4> ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0205.Ivo1  ( .en(GND), .in(\ILAB0606.ILE0205.net2656 ), .out(\ILAB0606.net15799 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0304.Iho1  ( .en(GND), .in(\ILAB0606.ILE0304.net2656 ), .out(\ILAB0606.net16132 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0304.Ivo1  ( .en(GND), .in(\ILAB0606.ILE0304.net2656 ), .out(\ILAB0606.net16114 ));
  inv_8_UCCLAB \ILAB0606.ILE0304.I666  ( .a(\ILAB0606.ILE0304.net0541 ), .x(\ILAB0606.net23576 ));
  inv_4_UCCLAB \ILAB0606.ILE0405.I713  ( .a(\ILAB0606.net23576 ), .x(\ILAB0606.ILE0405.net01342 ));
  inv_4_UCCLAB \ILAB0606.ILE0403.I715  ( .a(\ILAB0606.net23576 ), .x(\ILAB0606.ILE0403.net01339 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0305.Iho3  ( .en(GND), .in(\ILAB0606.ILE0305.net2656 ), .out(\ILAB0606.net23334 ));
  inv_8_UCCLAB \ILAB0606.ILE0405.I666  ( .a(\ILAB0606.ILE0405.net0541 ), .x(\ILAB0606.net15566 ));
  inv_4_UCCLAB \ILAB0606.ILE0506.I715  ( .a(\ILAB0606.net15566 ), .x(\ILAB0606.ILE0506.net01339 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0506.Ivi7  ( .en(GND), .in(\ILAB0606.ILE0506.net2656 ), .out(\net15022<5> ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0404.Ihi5  ( .en(GND), .in(\ILAB0606.ILE0404.net2656 ), .out(\ILAB0606.net26213 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0403.Ihi5  ( .en(GND), .in(\ILAB0606.ILE0403.net2656 ), .out(\ILAB0606.net20723 ));
  inv_8_UCCLAB \ILAB0606.ILE0403.I666  ( .a(\ILAB0606.ILE0403.net0541 ), .x(\ILAB0606.net26231 ));
  inv_4_UCCLAB \ILAB0606.ILE0502.I715  ( .a(\ILAB0606.net26231 ), .x(\ILAB0606.ILE0502.net01339 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0403.Ihi6  ( .en(GND), .in(\ILAB0606.ILE0403.net2656 ), .out(\net14051<6> ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0403.Ivo2  ( .en(GND), .in(\ILAB0606.ILE0403.net2656 ), .out(\ILAB0606.net17687 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0502.Ivi7  ( .en(GND), .in(\ILAB0606.ILE0502.net2656 ), .out(\net15022<1> ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0503.Iho1  ( .en(GND), .in(\ILAB0606.ILE0503.net2656 ), .out(\ILAB0606.net20137 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0505.Ihi7  ( .en(GND), .in(\ILAB0606.ILE0505.net2656 ), .out(\ILAB0606.net20632 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0501.Ihi5  ( .en(GND), .in(\ILAB0606.ILE0501.net2656 ), .out(\net14047<2> ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0501.Ihi6  ( .en(GND), .in(\ILAB0606.ILE0501.net2656 ), .out(\net14047<1> ));
  inv_8_UCCLAB \ILAB0606.ILE0501.I666  ( .a(\ILAB0606.ILE0501.net0541 ), .x(\net13981<0> ));
  inv_4_UCCLAB \ILAB0605.ILE0616.I713  ( .a(\net13981<0> ), .x(\ILAB0605.ILE0616.net01342 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE0501.Ihi7  ( .en(GND), .in(\ILAB0606.ILE0501.net2656 ), .out(\net14047<0> ));
  inv_8_UCCLAB \ILAB0606.ILE0401.I666  ( .a(\ILAB0606.ILE0401.net0541 ), .x(\net13982<0> ));
  inv_4_UCCLAB \ILAB0605.ILE0516.I715  ( .a(\net13982<0> ), .x(\ILAB0605.ILE0516.net01339 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0516.Ihi7  ( .en(GND), .in(\ILAB0605.ILE0516.net2656 ), .out(\ILAB0605.net19057 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0615.Iho3  ( .en(GND), .in(\ILAB0605.ILE0615.net2656 ), .out(\ILAB0605.net23964 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0616.Iho3  ( .en(GND), .in(\ILAB0605.ILE0616.net2656 ), .out(\net14043<4> ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0614.Ivi7  ( .en(GND), .in(\ILAB0605.ILE0614.net2656 ), .out(\ILAB0605.net22144 ));
  inv_8_UCCLAB \ILAB0605.ILE0614.I666  ( .a(\ILAB0605.ILE0614.net0541 ), .x(\ILAB0605.net19346 ));
  inv_4_UCCLAB \ILAB0605.ILE0513.I712  ( .a(\ILAB0605.net19346 ), .x(\ILAB0605.ILE0513.net0562 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0614.Ihi6  ( .en(GND), .in(\ILAB0605.ILE0614.net2656 ), .out(\ILAB0605.net21442 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0611.Ihi7  ( .en(GND), .in(\ILAB0605.net21442 ), .out(\ILAB0605.net17077 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0410.Ihi7  ( .en(GND), .in(\ILAB0605.net22144 ), .out(\ILAB0605.net18112 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0514.Ihi7  ( .en(GND), .in(\ILAB0605.ILE0514.net2656 ), .out(\ILAB0605.net23917 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0513.Ivo1  ( .en(GND), .in(\ILAB0605.ILE0513.net2656 ), .out(\ILAB0605.net25519 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0411.Ihi7  ( .en(GND), .in(\ILAB0605.ILE0411.net2656 ), .out(\ILAB0605.net16672 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0410.Ivo1  ( .en(GND), .in(\ILAB0605.ILE0410.net2656 ), .out(\ILAB0605.net23629 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0611.Iho3  ( .en(GND), .in(\ILAB0605.ILE0611.net2656 ), .out(\ILAB0605.net21444 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0512.Ivo1  ( .en(GND), .in(\ILAB0605.ILE0512.net2656 ), .out(\ILAB0605.net18949 ));
  inv_8_UCCLAB \ILAB0605.ILE0612.I666  ( .a(\ILAB0605.ILE0612.net0541 ), .x(\ILAB0605.net21461 ));
  inv_4_UCCLAB \ILAB0605.ILE0711.I714  ( .a(\ILAB0605.net21461 ), .x(\ILAB0605.ILE0711.net01345 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0412.Ivi7  ( .en(GND), .in(\ILAB0605.ILE0412.net2656 ), .out(\net14018<6> ));
  inv_8_UCCLAB \ILAB0605.ILE0413.I666  ( .a(\ILAB0605.ILE0413.net0541 ), .x(\ILAB0605.net19031 ));
  inv_4_UCCLAB \ILAB0605.ILE0312.I710  ( .a(\ILAB0605.net19031 ), .x(\ILAB0605.ILE0312.net0558 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0413.Ivi7  ( .en(GND), .in(\ILAB0605.ILE0413.net2656 ), .out(\net14014<6> ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0312.Iho3  ( .en(GND), .in(\ILAB0605.ILE0312.net2656 ), .out(\ILAB0605.net24909 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0211.Ivo1  ( .en(GND), .in(\ILAB0605.ILE0211.net2656 ), .out(\ILAB0605.net21469 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0311.Ihi7  ( .en(GND), .in(\ILAB0605.ILE0311.net2656 ), .out(\ILAB0605.net25852 ));
  inv_8_UCCLAB \ILAB0605.ILE0213.I666  ( .a(\ILAB0605.ILE0213.net0541 ), .x(\ILAB0605.net22316 ));
  inv_4_UCCLAB \ILAB0605.ILE0112.I712  ( .a(\ILAB0605.net22316 ), .x(\ILAB0605.ILE0112.net0562 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0212.Ivi7  ( .en(GND), .in(\ILAB0605.ILE0212.net2656 ), .out(\net14018<1> ));
  inv_8_UCCLAB \ILAB0605.ILE0212.I666  ( .a(\ILAB0605.ILE0212.net0541 ), .x(\ILAB0605.net23306 ));
  inv_4_UCCLAB \ILAB0605.ILE0111.I711  ( .a(\ILAB0605.net23306 ), .x(\ILAB0605.ILE0111.net0560 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0112.Iho3  ( .en(GND), .in(\ILAB0605.ILE0112.net2656 ), .out(\ILAB0605.net21894 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0111.Ihi7  ( .en(GND), .in(\ILAB0605.ILE0111.net2656 ), .out(\ILAB0605.net16807 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0110.Ivi7  ( .en(GND), .in(\ILAB0605.ILE0110.net2656 ), .out(\net14026<0> ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1612.Ivi7  ( .en(GND), .in(\ILAB0505.ILE1612.net2656 ), .out(\net13659<3> ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1611.Ivi7  ( .en(GND), .in(\ILAB0505.ILE1611.net2656 ), .out(\net13659<2> ));
  inv_8_UCCLAB \ILAB0505.ILE1611.I666  ( .a(\ILAB0505.ILE1611.net0541 ), .x(\ILAB0505.net24386 ));
  buftd4_UCCLAB \ILAB0505.I196  ( .a(\ILAB0505.net24386 ), .en(VDD), .x(\ILAB0505.net015234 ));
  mux2p_2_UCCLAB \ILAB0505.I5605.I0  ( .d0(GND), .d1(\ILAB0505.net015234 ), .s0(VDD), .x(\ILAB0505.I5605.net29 ));
  invd16_seth_UCCLAB \ILAB0505.I5605.I1  ( .a(\ILAB0505.I5605.net29 ), .c(VDD), .x(\ILAB0505.Clk_int<3> ));
  mux2d1i_1_P_UCCLAB \ILAB0505.I5366.I81  ( .d0(\ILAB0505.Clk_int<3> ), .d1i(GND), .sl0(GND), .x(\ILAB0505.I5366.net0102 ));
  invd52_UCCLAB \ILAB0505.I5366.I77  ( .a(\ILAB0505.I5366.net0102 ), .x(\ILAB0505.net15299<0> ));
  invd32_UCCLAB \ILAB0505.I5591.I0  ( .a(\ILAB0505.net15299<0> ), .x(\ILAB0505.Clk_LAB<3> ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1512.Ihi7  ( .en(GND), .in(\ILAB0505.ILE1512.net2656 ), .out(\ILAB0505.net19552 ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1411.Iho3  ( .en(GND), .in(\ILAB0505.ILE1411.net2656 ), .out(\ILAB0505.net20409 ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1412.Ivi7  ( .en(GND), .in(\ILAB0505.ILE1412.net2656 ), .out(\ILAB0505.net19399 ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1413.Ivi7  ( .en(GND), .in(\ILAB0505.ILE1413.net2656 ), .out(\ILAB0505.net18364 ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1513.Ivi7  ( .en(GND), .in(\ILAB0505.ILE1513.net2656 ), .out(\ILAB0505.net19219 ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1513.Iho1  ( .en(GND), .in(\ILAB0505.ILE1513.net2656 ), .out(\net13705<0> ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1513.Ivi5  ( .en(GND), .in(\ILAB0505.ILE1513.net2656 ), .out(\ILAB0505.net19217 ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1316.Iho2  ( .en(GND), .in(\ILAB0505.net19217 ), .out(\net13713<5> ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1313.Iho3  ( .en(GND), .in(\ILAB0505.ILE1313.net2656 ), .out(\ILAB0505.net20994 ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1416.Ivi7  ( .en(GND), .in(\ILAB0505.ILE1416.net2656 ), .out(\ILAB0505.net17914 ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1316.Ihi5  ( .en(GND), .in(\ILAB0505.ILE1316.net2656 ), .out(\ILAB0505.net23243 ));
  inv_8_UCCLAB \ILAB0505.ILE1316.I666  ( .a(\ILAB0505.ILE1316.net0541 ), .x(\net13671<1> ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1316.Ivi5  ( .en(GND), .in(\ILAB0505.ILE1316.net2656 ), .out(\ILAB0505.net20972 ));
  inv_4_UCCLAB \ILAB0505.ILE1215.I711  ( .a(\net13671<1> ), .x(\ILAB0505.ILE1215.net0560 ));
  inv_4_UCCLAB \ILAB0506.ILE1201.I711  ( .a(\net13671<1> ), .x(\ILAB0506.ILE1201.net0560 ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1216.Ihi7  ( .en(GND), .in(\ILAB0505.ILE1216.net2656 ), .out(\ILAB0505.net21352 ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1315.Ivi7  ( .en(GND), .in(\ILAB0505.ILE1315.net2656 ), .out(\ILAB0505.net24304 ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1215.Ivi7  ( .en(GND), .in(\ILAB0505.ILE1215.net2656 ), .out(\ILAB0505.net24439 ));
  inv_8_UCCLAB \ILAB0506.ILE1201.I666  ( .a(\ILAB0506.ILE1201.net0541 ), .x(\net13672<0> ));
  inv_4_UCCLAB \ILAB0506.ILE1302.I713  ( .a(\net13672<0> ), .x(\ILAB0506.ILE1302.net01342 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1501.Iho1  ( .en(GND), .in(\ILAB0506.ILE1501.net2656 ), .out(\ILAB0506.net20857 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1401.Iho3  ( .en(GND), .in(\ILAB0506.ILE1401.net2656 ), .out(\ILAB0506.net20814 ));
  inv_8_UCCLAB \ILAB0506.ILE1401.I666  ( .a(\ILAB0506.ILE1401.net0541 ), .x(\net13670<0> ));
  inv_4_UCCLAB \ILAB0506.ILE1302.I710  ( .a(\net13670<0> ), .x(\ILAB0506.ILE1302.net0558 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1302.Ivi7  ( .en(GND), .in(\ILAB0506.ILE1302.net2656 ), .out(\ILAB0506.net26554 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1403.Ihi7  ( .en(GND), .in(\ILAB0506.ILE1403.net2656 ), .out(\net13709<3> ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1402.Iho1  ( .en(GND), .in(\ILAB0506.ILE1402.net2656 ), .out(\ILAB0506.net26302 ));
  inv_8_UCCLAB \ILAB0506.ILE1504.I666  ( .a(\ILAB0506.ILE1504.net0541 ), .x(\ILAB0506.net17726 ));
  inv_4_UCCLAB \ILAB0506.ILE1603.I714  ( .a(\ILAB0506.net17726 ), .x(\ILAB0506.ILE1603.net01345 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1503.Ihi7  ( .en(GND), .in(\ILAB0506.ILE1503.net2656 ), .out(\net13705<3> ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1503.Ihi6  ( .en(GND), .in(\ILAB0506.ILE1503.net2656 ), .out(\net13705<6> ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1503.Ivi6  ( .en(GND), .in(\ILAB0506.ILE1503.net2656 ), .out(\ILAB0506.net15484 ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1516.Ihi7  ( .en(GND), .in(\net13705<6> ), .out(\ILAB0505.net19642 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1603.Iho3  ( .en(GND), .in(\ILAB0506.ILE1603.net2656 ), .out(\ILAB0506.net15459 ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1615.Ivi7  ( .en(GND), .in(\ILAB0505.ILE1615.net2656 ), .out(\net13659<6> ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1515.Ivi7  ( .en(GND), .in(\ILAB0505.ILE1515.net2656 ), .out(\ILAB0505.net22819 ));
  inv_8_UCCLAB \ILAB0505.ILE1516.I666  ( .a(\ILAB0505.ILE1516.net0541 ), .x(\net13669<1> ));
  inv_4_UCCLAB \ILAB0506.ILE1601.I713  ( .a(\net13669<1> ), .x(\ILAB0506.ILE1601.net01342 ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1616.Ivi6  ( .en(GND), .in(\ILAB0505.ILE1616.net2656 ), .out(\net14002<0> ));
  sw_b_v2_inv_UCCLAB \ILAB0505.ILE1616.Iho2  ( .en(GND), .in(\ILAB0505.ILE1616.net2656 ), .out(\net13701<5> ));
  inv_8_UCCLAB \ILAB0506.ILE1601.I666  ( .a(\ILAB0506.ILE1601.net0541 ), .x(\net13668<0> ));
  buftd4_UCCLAB \ILAB0506.I236  ( .a(\net13668<0> ), .en(VDD), .x(\ILAB0506.net027166 ));
  mux2p_2_UCCLAB \ILAB0506.I5605.I4  ( .d0(\ILAB0506.net027166 ), .d1(GND), .s0(GND), .x(\ILAB0506.I5605.net25 ));
  invd16_seth_UCCLAB \ILAB0506.I5605.I5  ( .a(\ILAB0506.I5605.net25 ), .c(VDD), .x(\ILAB0506.Clk_int<1> ));
  mux2d1i_1_P_UCCLAB \ILAB0506.I5366.I79  ( .d0(\ILAB0506.Clk_int<1> ), .d1i(GND), .sl0(GND), .x(\ILAB0506.I5366.net0110 ));
  invd52_UCCLAB \ILAB0506.I5366.I75  ( .a(\ILAB0506.I5366.net0110 ), .x(\ILAB0506.net15299<2> ));
  invd32_UCCLAB \ILAB0506.I5591.I2  ( .a(\ILAB0506.net15299<2> ), .x(\ILAB0506.Clk_LAB<1> ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0116.Ihi7  ( .en(GND), .in(\ILAB0605.ILE0116.net2656 ), .out(\ILAB0605.net21892 ));
  sw_b_v2_inv_UCCLAB \ILAB0605.ILE0115.Ivo3  ( .en(GND), .in(\ILAB0605.ILE0115.net2656 ), .out(\ILAB0605.net24615 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1112.Iho3  ( .en(GND), .in(\ILAB0506.ILE1112.net2656 ), .out(\ILAB0506.net21759 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1014.Ihi7  ( .en(GND), .in(\ILAB0506.ILE1014.net2656 ), .out(\ILAB0506.net24862 ));
  inv_8_UCCLAB \ILAB0506.ILE1014.I666  ( .a(\ILAB0506.ILE1014.net0541 ), .x(\ILAB0506.net21416 ));
  inv_4_UCCLAB \ILAB0506.ILE1113.I715  ( .a(\ILAB0506.net21416 ), .x(\ILAB0506.ILE1113.net01339 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1113.Iho3  ( .en(GND), .in(\ILAB0506.ILE1113.net2656 ), .out(\ILAB0506.net21534 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1013.Ivi7  ( .en(GND), .in(\ILAB0506.ILE1013.net2656 ), .out(\ILAB0506.net21424 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1012.Ivi7  ( .en(GND), .in(\ILAB0506.ILE1012.net2656 ), .out(\ILAB0506.net21694 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE1012.Ivi5  ( .en(GND), .in(\ILAB0506.ILE1012.net2656 ), .out(\ILAB0506.net21692 ));
  inv_8_UCCLAB \ILAB0506.ILE1012.I666  ( .a(\ILAB0506.ILE1012.net0541 ), .x(\ILAB0506.net22676 ));
  inv_4_UCCLAB \ILAB0506.ILE0913.I712  ( .a(\ILAB0506.net22676 ), .x(\ILAB0506.ILE0913.net0562 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE0915.Ihi5  ( .en(GND), .in(\ILAB0506.ILE0915.net2656 ), .out(\ILAB0506.net25493 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE0913.Ihi7  ( .en(GND), .in(\ILAB0506.ILE0913.net2656 ), .out(\ILAB0506.net25312 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE0813.Ivi7  ( .en(GND), .in(\ILAB0506.ILE0813.net2656 ), .out(\ILAB0506.net22549 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE0914.Ivi6  ( .en(GND), .in(\ILAB0506.ILE0914.net2656 ), .out(\ILAB0506.net23494 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE0713.Iho3  ( .en(GND), .in(\ILAB0506.ILE0713.net2656 ), .out(\ILAB0506.net19959 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE0712.Ivi7  ( .en(GND), .in(\ILAB0506.ILE0712.net2656 ), .out(\ILAB0506.net19939 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE0613.Ihi5  ( .en(GND), .in(\ILAB0506.ILE0613.net2656 ), .out(\ILAB0506.net21443 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE0613.Ivi7  ( .en(GND), .in(\ILAB0506.ILE0613.net2656 ), .out(\ILAB0506.net19354 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE0612.Ihi5  ( .en(GND), .in(\ILAB0506.ILE0612.net2656 ), .out(\ILAB0506.net24098 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE0311.Ivo1  ( .en(GND), .in(\ILAB0506.ILE0311.net2656 ), .out(\ILAB0506.net21514 ));
  inv_8_UCCLAB \ILAB0506.ILE0312.I666  ( .a(\ILAB0506.ILE0312.net0541 ), .x(\ILAB0506.net23396 ));
  inv_4_UCCLAB \ILAB0506.ILE0411.I715  ( .a(\ILAB0506.net23396 ), .x(\ILAB0506.ILE0411.net01339 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE0312.Ivi6  ( .en(GND), .in(\ILAB0506.ILE0312.net2656 ), .out(\net14773<6> ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE0411.Ivo1  ( .en(GND), .in(\ILAB0506.ILE0411.net2656 ), .out(\ILAB0506.net18499 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE0412.Iho3  ( .en(GND), .in(\ILAB0506.ILE0412.net2656 ), .out(\ILAB0506.net19014 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE0313.Iho1  ( .en(GND), .in(\ILAB0506.ILE0313.net2656 ), .out(\net14810<0> ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE0313.Ivo1  ( .en(GND), .in(\ILAB0506.ILE0313.net2656 ), .out(\ILAB0506.net19984 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE0313.Iho2  ( .en(GND), .in(\ILAB0506.ILE0313.net2656 ), .out(\ILAB0506.net23153 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE0315.Iho3  ( .en(GND), .in(\ILAB0506.net23153 ), .out(\ILAB0506.net24819 ));
  inv_8_UCCLAB \ILAB0506.ILE0413.I666  ( .a(\ILAB0506.ILE0413.net0541 ), .x(\ILAB0506.net19031 ));
  inv_4_UCCLAB \ILAB0506.ILE0512.I714  ( .a(\ILAB0506.net19031 ), .x(\ILAB0506.ILE0512.net01345 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE0314.Ivo1  ( .en(GND), .in(\ILAB0506.ILE0314.net2656 ), .out(\ILAB0506.net22414 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE0415.Ivo1  ( .en(GND), .in(\ILAB0506.ILE0415.net2656 ), .out(\ILAB0506.net22099 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE0415.Ihi5  ( .en(GND), .in(\ILAB0506.ILE0415.net2656 ), .out(\ILAB0506.net26078 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE0414.Ivo1  ( .en(GND), .in(\ILAB0506.ILE0414.net2656 ), .out(\ILAB0506.net18904 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE0515.Ivo1  ( .en(GND), .in(\ILAB0506.ILE0515.net2656 ), .out(\ILAB0506.net22189 ));
  sw_b_v2_inv_UCCLAB \ILAB0506.ILE0615.Ihi7  ( .en(GND), .in(\ILAB0506.ILE0615.net2656 ), .out(\ILAB0506.net21442 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1309.Ivi7  ( .en(GND), .in(\ILAB0606.ILE1309.net2656 ), .out(\ILAB0606.net16249 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1309.Iho1  ( .en(GND), .in(\ILAB0606.ILE1309.net2656 ), .out(\ILAB0606.net16222 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1309.Ivi6  ( .en(GND), .in(\ILAB0606.ILE1309.net2656 ), .out(\ILAB0606.net18094 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1309.Ivo2  ( .en(GND), .in(\ILAB0606.ILE1309.net2656 ), .out(\ILAB0606.net18047 ));
  inv_8_UCCLAB \ILAB0606.ILE1309.I666  ( .a(\ILAB0606.ILE1309.net0541 ), .x(\ILAB0606.net21866 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1209.Ivo2  ( .en(GND), .in(\ILAB0606.net16249 ), .out(\ILAB0606.net18092 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1409.Ivo1  ( .en(GND), .in(\ILAB0606.net18094 ), .out(\net14936<1> ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1509.Ivo3  ( .en(GND), .in(\ILAB0606.net18047 ), .out(\ILAB0606.net16020 ));
  inv_4_UCCLAB \ILAB0606.ILE1410.I714  ( .a(\ILAB0606.net21866 ), .x(\ILAB0606.ILE1410.net01345 ));
  inv_4_UCCLAB \ILAB0606.ILE1410.I715  ( .a(\ILAB0606.net21866 ), .x(\ILAB0606.ILE1410.net01339 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1412.Iho2  ( .en(GND), .in(\net14936<1> ), .out(\ILAB0606.net19373 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1312.Iho2  ( .en(GND), .in(\ILAB0606.net16222 ), .out(\ILAB0606.net21218 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1512.Iho2  ( .en(GND), .in(\ILAB0606.net16020 ), .out(\ILAB0606.net19643 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1209.Ivi5  ( .en(GND), .in(\ILAB0606.ILE1209.net2656 ), .out(\ILAB0606.net16292 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1109.Ivo1  ( .en(GND), .in(\ILAB0606.ILE1109.net2656 ), .out(\ILAB0606.net18049 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1210.Ivo2  ( .en(GND), .in(\ILAB0606.ILE1210.net2656 ), .out(\ILAB0606.net24032 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1410.Ivo3  ( .en(GND), .in(\ILAB0606.net24032 ), .out(\ILAB0606.net24075 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1210.Iho2  ( .en(GND), .in(\ILAB0606.ILE1210.net2656 ), .out(\ILAB0606.net24728 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1212.Iho3  ( .en(GND), .in(\ILAB0606.net24728 ), .out(\ILAB0606.net21354 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1210.Iho3  ( .en(GND), .in(\ILAB0606.ILE1210.net2656 ), .out(\ILAB0606.net24729 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1311.Ivo1  ( .en(GND), .in(\ILAB0606.net24729 ), .out(\net14928<0> ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1413.Iho2  ( .en(GND), .in(\ILAB0606.net24075 ), .out(\ILAB0606.net18338 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1310.Iho3  ( .en(GND), .in(\ILAB0606.ILE1310.net2656 ), .out(\ILAB0606.net24684 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1310.Iho1  ( .en(GND), .in(\ILAB0606.ILE1310.net2656 ), .out(\ILAB0606.net24682 ));
  inv_8_UCCLAB \ILAB0606.ILE1310.I666  ( .a(\ILAB0606.ILE1310.net0541 ), .x(\ILAB0606.net16241 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1313.Iho2  ( .en(GND), .in(\ILAB0606.net24682 ), .out(\ILAB0606.net20993 ));
  inv_4_UCCLAB \ILAB0606.ILE1411.I715  ( .a(\ILAB0606.net16241 ), .x(\ILAB0606.ILE1411.net01339 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1310.Ivo1  ( .en(GND), .in(\ILAB0606.ILE1310.net2656 ), .out(\net14932<0> ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1310.Ivo2  ( .en(GND), .in(\ILAB0606.ILE1310.net2656 ), .out(\ILAB0606.net24077 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1610.Ivo2  ( .en(GND), .in(\net14932<0> ), .out(\net14932<5> ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1510.Ivo3  ( .en(GND), .in(\ILAB0606.net24077 ), .out(\ILAB0606.net24390 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1312.Iho3  ( .en(GND), .in(\ILAB0606.ILE1312.net2656 ), .out(\ILAB0606.net21219 ));
  inv_8_UCCLAB \ILAB0606.ILE1312.I666  ( .a(\ILAB0606.ILE1312.net0541 ), .x(\ILAB0606.net22226 ));
  inv_4_UCCLAB \ILAB0606.ILE1213.I710  ( .a(\ILAB0606.net22226 ), .x(\ILAB0606.ILE1213.net0558 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1312.Ivi5  ( .en(GND), .in(\ILAB0606.ILE1312.net2656 ), .out(\ILAB0606.net21242 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1114.Ivo1  ( .en(GND), .in(\ILAB0606.ILE1114.net2656 ), .out(\ILAB0606.net22054 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1114.Ihi6  ( .en(GND), .in(\ILAB0606.ILE1114.net2656 ), .out(\ILAB0606.net23017 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1114.Ihi5  ( .en(GND), .in(\ILAB0606.ILE1114.net2656 ), .out(\ILAB0606.net21758 ));
  inv_8_UCCLAB \ILAB0606.ILE1114.I666  ( .a(\ILAB0606.ILE1114.net0541 ), .x(\ILAB0606.net21551 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1414.Ivo2  ( .en(GND), .in(\ILAB0606.net22054 ), .out(\ILAB0606.net22772 ));
  inv_4_UCCLAB \ILAB0606.ILE1213.I714  ( .a(\ILAB0606.net21551 ), .x(\ILAB0606.ILE1213.net01345 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1614.Ivo3  ( .en(GND), .in(\ILAB0606.net22772 ), .out(\net14916<4> ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1213.Iho2  ( .en(GND), .in(\ILAB0606.net22054 ), .out(\ILAB0606.net21083 ));
  inv_8_UCCLAB \ILAB0606.ILE1314.I666  ( .a(\ILAB0606.net22054 ), .x(\ILAB0606.net21011 ));
  inv_8_UCCLAB \ILAB0606.ILE1212.I666  ( .a(\ILAB0606.ILE1212.net0541 ), .x(\ILAB0606.net22586 ));
  inv_4_UCCLAB \ILAB0606.ILE1111.I712  ( .a(\ILAB0606.net22586 ), .x(\ILAB0606.ILE1111.net0562 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1410.Ivo2  ( .en(GND), .in(\ILAB0606.ILE1410.net2656 ), .out(\ILAB0606.net24392 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1610.Ivo3  ( .en(GND), .in(\ILAB0606.net24392 ), .out(\net14932<4> ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1410.Ivi7  ( .en(GND), .in(\ILAB0606.ILE1410.net2656 ), .out(\ILAB0606.net24034 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1111.Ihi5  ( .en(GND), .in(\ILAB0606.ILE1111.net2656 ), .out(\ILAB0606.net16358 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1110.Ivo1  ( .en(GND), .in(\ILAB0606.ILE1110.net2656 ), .out(\ILAB0606.net24079 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1211.Ivo1  ( .en(GND), .in(\ILAB0606.ILE1211.net2656 ), .out(\net15018<2> ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1412.Ivi7  ( .en(GND), .in(\ILAB0606.ILE1412.net2656 ), .out(\ILAB0606.net19399 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1412.Iho1  ( .en(GND), .in(\ILAB0606.ILE1412.net2656 ), .out(\ILAB0606.net19372 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1412.Ivi5  ( .en(GND), .in(\ILAB0606.ILE1412.net2656 ), .out(\ILAB0606.net19397 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1415.Iho2  ( .en(GND), .in(\ILAB0606.net19372 ), .out(\net15068<2> ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1112.Ihi7  ( .en(GND), .in(\ILAB0606.ILE1112.net2656 ), .out(\ILAB0606.net24772 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1111.Iho2  ( .en(GND), .in(\ILAB0606.net24772 ), .out(\ILAB0606.net23018 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1311.Ihi7  ( .en(GND), .in(\ILAB0606.ILE1311.net2656 ), .out(\ILAB0606.net17122 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1213.Ivi7  ( .en(GND), .in(\ILAB0606.ILE1213.net2656 ), .out(\ILAB0606.net21109 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1411.Ivo1  ( .en(GND), .in(\ILAB0606.ILE1411.net2656 ), .out(\net14928<1> ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1214.Ivi7  ( .en(GND), .in(\ILAB0606.ILE1214.net2656 ), .out(\ILAB0606.net23449 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1014.Ihi7  ( .en(GND), .in(\ILAB0606.ILE1014.net2656 ), .out(\ILAB0606.net24862 ));
  inv_8_UCCLAB \ILAB0606.ILE1013.I666  ( .a(\ILAB0606.ILE1013.net0541 ), .x(\ILAB0606.net21686 ));
  inv_4_UCCLAB \ILAB0606.ILE1114.I714  ( .a(\ILAB0606.net21686 ), .x(\ILAB0606.ILE1114.net01345 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1413.Iho1  ( .en(GND), .in(\ILAB0606.ILE1413.net2656 ), .out(\net15068<0> ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1513.Iho1  ( .en(GND), .in(\ILAB0606.ILE1513.net2656 ), .out(\net15064<0> ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1414.Ivo1  ( .en(GND), .in(\ILAB0606.ILE1414.net2656 ), .out(\net14916<1> ));
  inv_8_UCCLAB \ILAB0606.ILE1414.I666  ( .a(\ILAB0606.ILE1414.net0541 ), .x(\ILAB0606.net18356 ));
  inv_4_UCCLAB \ILAB0606.ILE1515.I714  ( .a(\ILAB0606.net18356 ), .x(\ILAB0606.ILE1515.net01345 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1511.Iho1  ( .en(GND), .in(\ILAB0606.ILE1511.net2656 ), .out(\ILAB0606.net21262 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1514.Ivo1  ( .en(GND), .in(\ILAB0606.ILE1514.net2656 ), .out(\net14916<3> ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1613.Ivo1  ( .en(GND), .in(\ILAB0606.ILE1613.net2656 ), .out(\net14920<6> ));
  inv_8_UCCLAB \ILAB0606.ILE1613.I666  ( .a(\ILAB0606.ILE1613.net0541 ), .x(\ILAB0606.net20111 ));
  buftd4_UCCLAB \ILAB0606.I189  ( .a(\ILAB0606.net20111 ), .en(VDD), .x(\ILAB0606.net27185 ));
  mux2p_2_UCCLAB \ILAB0606.I5605.I7  ( .d0(GND), .d1(\ILAB0606.net27185 ), .s0(VDD), .x(\ILAB0606.I5605.net21 ));
  invd16_seth_UCCLAB \ILAB0606.I5605.I6  ( .a(\ILAB0606.I5605.net21 ), .c(VDD), .x(\ILAB0606.Clk_int<0> ));
  mux2p_2_UCCLAB \ILAB0606.I5366.I82  ( .d0(\ILAB0606.Clk_int<0> ), .d1(GND), .s0(GND), .x(\ILAB0606.I5366.net0119 ));
  invtd56_clk_UCCLAB \ILAB0606.I5366.I6  ( .a(\ILAB0606.I5366.net0119 ), .en(VDD), .x(\net10229<1> ));
  invtd56_UCCLAB \I3692.I4  ( .a(\net10229<1> ), .en(VDD), .x(\net10255<1> ));
  mux2p_2_UCCLAB \I3686.I2  ( .d0(GND), .d1(\net10255<1> ), .s0(VDD), .x(\I3686.net35 ));
  invtd56_pd_clk_UCCLAB \I3686.I9  ( .a(\I3686.net35 ), .en(VDD), .x(\net10252<3> ));
  invtd56_pd_clk_UCCLAB \I3637.I4  ( .a(\net10252<3> ), .en(VDD), .x(\net20148<3> ));
  nand2_1_UCCLAB \ILAB0706.I5366.I0  ( .a(VDD), .b(\net20148<3> ), .x(\ILAB0706.I5366.net64 ));
  mux2d1i_1_P_UCCLAB \ILAB0706.I5366.I78  ( .d0(GND), .d1i(\ILAB0706.I5366.net64 ), .sl0(VDD), .x(\ILAB0706.I5366.net0114 ));
  invd52_UCCLAB \ILAB0706.I5366.I74  ( .a(\ILAB0706.I5366.net0114 ), .x(\ILAB0706.net15299<3> ));
  invd32_UCCLAB \ILAB0706.I5591.I3  ( .a(\ILAB0706.net15299<3> ), .x(\ILAB0706.Clk_LAB<0> ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1512.Ivo2  ( .en(GND), .in(\ILAB0606.ILE1512.net2656 ), .out(\net14924<2> ));
  sw_b_v2_inv_UCCLAB \ILAB0706.ILE0112.Ivo3  ( .en(GND), .in(\net14924<2> ), .out(\ILAB0706.net22320 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1612.Iho1  ( .en(GND), .in(\ILAB0606.ILE1612.net2656 ), .out(\ILAB0606.net20092 ));
  sw_b_v2_inv_UCCLAB \ILAB0606.ILE1614.Ivo1  ( .en(GND), .in(\ILAB0606.ILE1614.net2656 ), .out(\net14916<6> ));
  inv_8_UCCLAB \ILAB0606.ILE1614.I666  ( .a(\ILAB0606.ILE1614.net0541 ), .x(\ILAB0606.net20066 ));
  buftd4_UCCLAB \ILAB0606.I183  ( .a(\ILAB0606.net20066 ), .en(VDD), .x(\ILAB0606.net27191 ));
  mux2p_2_UCCLAB \ILAB0606.I5605.I4  ( .d0(GND), .d1(\ILAB0606.net27191 ), .s0(VDD), .x(\ILAB0606.I5605.net25 ));
  invd16_seth_UCCLAB \ILAB0606.I5605.I5  ( .a(\ILAB0606.I5605.net25 ), .c(VDD), .x(\ILAB0606.Clk_int<1> ));
  mux2p_2_UCCLAB \ILAB0606.I5366.I83  ( .d0(\ILAB0606.Clk_int<1> ), .d1(GND), .s0(GND), .x(\ILAB0606.I5366.net0122 ));
  invtd56_clk_UCCLAB \ILAB0606.I5366.I8  ( .a(\ILAB0606.I5366.net0122 ), .en(VDD), .x(\net10229<0> ));
  invtd56_UCCLAB \I3692.I3  ( .a(\net10229<0> ), .en(VDD), .x(\net10255<0> ));
  mux2p_2_UCCLAB \I3686.I3  ( .d0(GND), .d1(\net10255<0> ), .s0(VDD), .x(\I3686.net39 ));
  invtd56_pd_clk_UCCLAB \I3686.I7  ( .a(\I3686.net39 ), .en(VDD), .x(\net10252<2> ));
  invtd56_pd_clk_UCCLAB \I3637.I3  ( .a(\net10252<2> ), .en(VDD), .x(\net20148<2> ));
  nand2_1_UCCLAB \ILAB0706.I5366.I71  ( .a(VDD), .b(\net20148<2> ), .x(\ILAB0706.I5366.net70 ));
  mux2d1i_1_P_UCCLAB \ILAB0706.I5366.I79  ( .d0(GND), .d1i(\ILAB0706.I5366.net70 ), .sl0(VDD), .x(\ILAB0706.I5366.net0110 ));
  invd52_UCCLAB \ILAB0706.I5366.I75  ( .a(\ILAB0706.I5366.net0110 ), .x(\ILAB0706.net15299<2> ));
  invd32_UCCLAB \ILAB0706.I5591.I2  ( .a(\ILAB0706.net15299<2> ), .x(\ILAB0706.Clk_LAB<1> ));
endmodule
///////////////////////////////////////////////////////
