//###########################################################
//##                                                         
//##   Created       X-CAD v2.74.68                               
//##   Date/Time     24.10.2024 / 11:12:11                                 
//##   Language      System Verilog                                      
//##                                                         
//###########################################################

module test();


endmodule
